VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_1
  CLASS BLOCK ;
  FOREIGN tt_um_test_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 43.460 BY 54.180 ;
  PIN Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.601000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END Out
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.245 10.640 14.245 41.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.295 10.640 22.295 41.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.345 10.640 30.345 41.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.395 10.640 38.395 41.740 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.315 38.395 19.315 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 24.790 38.395 26.790 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 32.265 38.395 34.265 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 39.740 38.395 41.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.545 10.640 10.545 41.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.595 10.640 18.595 41.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.645 10.640 26.645 41.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.695 10.640 34.695 41.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 13.615 37.960 15.615 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 21.090 37.960 23.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 28.565 37.960 30.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 36.040 37.960 38.040 ;
    END
  END VPWR
  PIN Vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END Vin
  PIN Vip
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END Vip
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END clk
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 37.910 40.990 ;
      LAYER li1 ;
        RECT 5.520 10.795 37.720 40.885 ;
      LAYER met1 ;
        RECT 4.210 10.640 38.395 41.040 ;
      LAYER met2 ;
        RECT 4.230 4.280 38.335 40.985 ;
        RECT 4.230 3.670 25.570 4.280 ;
        RECT 26.410 3.670 38.335 4.280 ;
      LAYER met3 ;
        RECT 3.990 28.240 38.385 40.965 ;
        RECT 4.400 26.840 38.385 28.240 ;
        RECT 3.990 24.840 38.385 26.840 ;
        RECT 4.400 23.440 38.385 24.840 ;
        RECT 3.990 10.715 38.385 23.440 ;
  END
END tt_um_test_1
END LIBRARY

