VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_brandonramos_opamp_ladder
  CLASS BLOCK ;
  FOREIGN tt_um_brandonramos_opamp_ladder ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  OBS
      LAYER pwell ;
        RECT 50.665 136.935 50.835 137.105 ;
        RECT 52.045 136.935 52.215 137.105 ;
        RECT 57.565 136.935 57.735 137.105 ;
        RECT 63.080 136.965 63.200 137.075 ;
        RECT 64.005 136.935 64.175 137.105 ;
        RECT 69.525 136.935 69.695 137.105 ;
        RECT 75.045 136.935 75.215 137.105 ;
        RECT 76.885 136.935 77.055 137.105 ;
        RECT 82.405 136.935 82.575 137.105 ;
        RECT 87.925 136.935 88.095 137.105 ;
        RECT 89.765 136.935 89.935 137.105 ;
        RECT 95.285 136.935 95.455 137.105 ;
        RECT 100.805 136.935 100.975 137.105 ;
        RECT 102.645 136.935 102.815 137.105 ;
        RECT 108.165 136.935 108.335 137.105 ;
        RECT 113.685 136.935 113.855 137.105 ;
        RECT 115.525 136.935 115.695 137.105 ;
        RECT 121.045 136.935 121.215 137.105 ;
        RECT 126.565 136.935 126.735 137.105 ;
        RECT 128.405 136.935 128.575 137.105 ;
        RECT 133.925 136.935 134.095 137.105 ;
        RECT 137.600 136.965 137.720 137.075 ;
        RECT 138.985 136.935 139.155 137.105 ;
        RECT 63.545 136.175 63.715 136.700 ;
        RECT 76.425 136.175 76.595 136.700 ;
        RECT 89.305 136.175 89.475 136.700 ;
        RECT 102.185 136.175 102.355 136.700 ;
        RECT 115.065 136.175 115.235 136.700 ;
        RECT 127.945 136.175 128.115 136.700 ;
      LAYER nwell ;
        RECT 50.330 132.885 139.490 135.715 ;
      LAYER pwell ;
        RECT 63.545 131.900 63.715 132.425 ;
        RECT 89.305 131.900 89.475 132.425 ;
        RECT 115.065 131.900 115.235 132.425 ;
        RECT 50.665 131.495 50.835 131.665 ;
        RECT 52.045 131.495 52.215 131.665 ;
        RECT 57.565 131.495 57.735 131.665 ;
        RECT 63.085 131.635 63.255 131.665 ;
        RECT 63.080 131.525 63.255 131.635 ;
        RECT 63.085 131.495 63.255 131.525 ;
        RECT 64.005 131.495 64.175 131.665 ;
        RECT 68.605 131.495 68.775 131.665 ;
        RECT 69.525 131.495 69.695 131.665 ;
        RECT 74.125 131.495 74.295 131.665 ;
        RECT 75.045 131.495 75.215 131.665 ;
        RECT 75.960 131.525 76.080 131.635 ;
        RECT 76.885 131.495 77.055 131.665 ;
        RECT 80.565 131.495 80.735 131.665 ;
        RECT 82.405 131.495 82.575 131.665 ;
        RECT 86.085 131.495 86.255 131.665 ;
        RECT 87.925 131.495 88.095 131.665 ;
        RECT 88.840 131.525 88.960 131.635 ;
        RECT 89.765 131.495 89.935 131.665 ;
        RECT 93.445 131.495 93.615 131.665 ;
        RECT 95.285 131.495 95.455 131.665 ;
        RECT 98.965 131.495 99.135 131.665 ;
        RECT 100.805 131.495 100.975 131.665 ;
        RECT 101.720 131.525 101.840 131.635 ;
        RECT 102.645 131.495 102.815 131.665 ;
        RECT 106.325 131.495 106.495 131.665 ;
        RECT 108.165 131.495 108.335 131.665 ;
        RECT 111.845 131.495 112.015 131.665 ;
        RECT 113.685 131.495 113.855 131.665 ;
        RECT 114.600 131.525 114.720 131.635 ;
        RECT 115.525 131.495 115.695 131.665 ;
        RECT 119.205 131.495 119.375 131.665 ;
        RECT 121.045 131.495 121.215 131.665 ;
        RECT 124.725 131.495 124.895 131.665 ;
        RECT 126.565 131.495 126.735 131.665 ;
        RECT 127.480 131.525 127.600 131.635 ;
        RECT 128.405 131.495 128.575 131.665 ;
        RECT 132.085 131.495 132.255 131.665 ;
        RECT 133.925 131.495 134.095 131.665 ;
        RECT 137.600 131.525 137.720 131.635 ;
        RECT 138.985 131.495 139.155 131.665 ;
        RECT 76.425 130.735 76.595 131.260 ;
        RECT 102.185 130.735 102.355 131.260 ;
        RECT 127.945 130.735 128.115 131.260 ;
      LAYER nwell ;
        RECT 50.330 127.445 139.490 130.275 ;
      LAYER pwell ;
        RECT 63.545 126.460 63.715 126.985 ;
        RECT 89.305 126.460 89.475 126.985 ;
        RECT 115.065 126.460 115.235 126.985 ;
        RECT 50.665 126.055 50.835 126.225 ;
        RECT 52.045 126.055 52.215 126.225 ;
        RECT 57.565 126.055 57.735 126.225 ;
        RECT 63.085 126.195 63.255 126.225 ;
        RECT 63.080 126.085 63.255 126.195 ;
        RECT 63.085 126.055 63.255 126.085 ;
        RECT 64.005 126.055 64.175 126.225 ;
        RECT 68.605 126.055 68.775 126.225 ;
        RECT 69.525 126.055 69.695 126.225 ;
        RECT 74.125 126.055 74.295 126.225 ;
        RECT 75.045 126.055 75.215 126.225 ;
        RECT 75.960 126.085 76.080 126.195 ;
        RECT 76.885 126.055 77.055 126.225 ;
        RECT 80.565 126.055 80.735 126.225 ;
        RECT 82.405 126.055 82.575 126.225 ;
        RECT 86.085 126.055 86.255 126.225 ;
        RECT 87.925 126.055 88.095 126.225 ;
        RECT 88.840 126.085 88.960 126.195 ;
        RECT 89.765 126.055 89.935 126.225 ;
        RECT 93.445 126.055 93.615 126.225 ;
        RECT 95.285 126.055 95.455 126.225 ;
        RECT 98.965 126.055 99.135 126.225 ;
        RECT 100.805 126.055 100.975 126.225 ;
        RECT 101.720 126.085 101.840 126.195 ;
        RECT 102.645 126.055 102.815 126.225 ;
        RECT 106.325 126.055 106.495 126.225 ;
        RECT 108.165 126.055 108.335 126.225 ;
        RECT 111.845 126.055 112.015 126.225 ;
        RECT 113.685 126.055 113.855 126.225 ;
        RECT 114.600 126.085 114.720 126.195 ;
        RECT 115.525 126.055 115.695 126.225 ;
        RECT 119.205 126.055 119.375 126.225 ;
        RECT 121.045 126.055 121.215 126.225 ;
        RECT 124.725 126.055 124.895 126.225 ;
        RECT 126.565 126.055 126.735 126.225 ;
        RECT 127.480 126.085 127.600 126.195 ;
        RECT 128.405 126.055 128.575 126.225 ;
        RECT 132.085 126.055 132.255 126.225 ;
        RECT 133.925 126.055 134.095 126.225 ;
        RECT 137.600 126.085 137.720 126.195 ;
        RECT 138.985 126.055 139.155 126.225 ;
        RECT 76.425 125.295 76.595 125.820 ;
        RECT 102.185 125.295 102.355 125.820 ;
        RECT 127.945 125.295 128.115 125.820 ;
      LAYER nwell ;
        RECT 50.330 122.005 139.490 124.835 ;
      LAYER pwell ;
        RECT 63.545 121.020 63.715 121.545 ;
        RECT 89.305 121.020 89.475 121.545 ;
        RECT 115.065 121.020 115.235 121.545 ;
        RECT 50.665 120.615 50.835 120.785 ;
        RECT 52.045 120.615 52.215 120.785 ;
        RECT 57.565 120.615 57.735 120.785 ;
        RECT 63.085 120.755 63.255 120.785 ;
        RECT 63.080 120.645 63.255 120.755 ;
        RECT 63.085 120.615 63.255 120.645 ;
        RECT 64.005 120.615 64.175 120.785 ;
        RECT 68.605 120.615 68.775 120.785 ;
        RECT 69.525 120.615 69.695 120.785 ;
        RECT 74.125 120.615 74.295 120.785 ;
        RECT 75.045 120.615 75.215 120.785 ;
        RECT 75.960 120.645 76.080 120.755 ;
        RECT 76.885 120.615 77.055 120.785 ;
        RECT 80.565 120.615 80.735 120.785 ;
        RECT 82.405 120.615 82.575 120.785 ;
        RECT 86.085 120.615 86.255 120.785 ;
        RECT 87.925 120.615 88.095 120.785 ;
        RECT 88.840 120.645 88.960 120.755 ;
        RECT 89.765 120.615 89.935 120.785 ;
        RECT 93.445 120.615 93.615 120.785 ;
        RECT 95.285 120.615 95.455 120.785 ;
        RECT 98.965 120.615 99.135 120.785 ;
        RECT 100.805 120.615 100.975 120.785 ;
        RECT 101.720 120.645 101.840 120.755 ;
        RECT 102.645 120.615 102.815 120.785 ;
        RECT 106.325 120.615 106.495 120.785 ;
        RECT 108.165 120.615 108.335 120.785 ;
        RECT 111.845 120.615 112.015 120.785 ;
        RECT 113.685 120.615 113.855 120.785 ;
        RECT 114.600 120.645 114.720 120.755 ;
        RECT 115.525 120.615 115.695 120.785 ;
        RECT 119.205 120.615 119.375 120.785 ;
        RECT 121.045 120.615 121.215 120.785 ;
        RECT 124.725 120.615 124.895 120.785 ;
        RECT 126.565 120.615 126.735 120.785 ;
        RECT 127.480 120.645 127.600 120.755 ;
        RECT 128.405 120.615 128.575 120.785 ;
        RECT 132.085 120.615 132.255 120.785 ;
        RECT 133.925 120.615 134.095 120.785 ;
        RECT 137.600 120.645 137.720 120.755 ;
        RECT 138.985 120.615 139.155 120.785 ;
        RECT 76.425 119.855 76.595 120.380 ;
        RECT 102.185 119.855 102.355 120.380 ;
        RECT 127.945 119.855 128.115 120.380 ;
      LAYER nwell ;
        RECT 50.330 116.565 139.490 119.395 ;
      LAYER pwell ;
        RECT 63.545 115.580 63.715 116.105 ;
        RECT 89.305 115.580 89.475 116.105 ;
        RECT 115.065 115.580 115.235 116.105 ;
        RECT 50.665 115.175 50.835 115.345 ;
        RECT 52.045 115.175 52.215 115.345 ;
        RECT 57.565 115.175 57.735 115.345 ;
        RECT 63.085 115.315 63.255 115.345 ;
        RECT 63.080 115.205 63.255 115.315 ;
        RECT 63.085 115.175 63.255 115.205 ;
        RECT 64.005 115.175 64.175 115.345 ;
        RECT 68.605 115.175 68.775 115.345 ;
        RECT 69.525 115.175 69.695 115.345 ;
        RECT 74.125 115.175 74.295 115.345 ;
        RECT 75.045 115.175 75.215 115.345 ;
        RECT 75.960 115.205 76.080 115.315 ;
        RECT 76.885 115.175 77.055 115.345 ;
        RECT 80.565 115.175 80.735 115.345 ;
        RECT 82.405 115.175 82.575 115.345 ;
        RECT 86.085 115.175 86.255 115.345 ;
        RECT 87.925 115.175 88.095 115.345 ;
        RECT 88.840 115.205 88.960 115.315 ;
        RECT 89.765 115.175 89.935 115.345 ;
        RECT 93.445 115.175 93.615 115.345 ;
        RECT 95.285 115.175 95.455 115.345 ;
        RECT 98.965 115.175 99.135 115.345 ;
        RECT 100.805 115.175 100.975 115.345 ;
        RECT 101.720 115.205 101.840 115.315 ;
        RECT 102.645 115.175 102.815 115.345 ;
        RECT 106.325 115.175 106.495 115.345 ;
        RECT 108.165 115.175 108.335 115.345 ;
        RECT 111.845 115.175 112.015 115.345 ;
        RECT 113.685 115.175 113.855 115.345 ;
        RECT 114.600 115.205 114.720 115.315 ;
        RECT 115.525 115.175 115.695 115.345 ;
        RECT 119.205 115.175 119.375 115.345 ;
        RECT 121.045 115.175 121.215 115.345 ;
        RECT 124.725 115.175 124.895 115.345 ;
        RECT 126.565 115.175 126.735 115.345 ;
        RECT 127.480 115.205 127.600 115.315 ;
        RECT 128.405 115.175 128.575 115.345 ;
        RECT 132.085 115.175 132.255 115.345 ;
        RECT 133.925 115.175 134.095 115.345 ;
        RECT 137.600 115.205 137.720 115.315 ;
        RECT 138.985 115.175 139.155 115.345 ;
        RECT 76.425 114.415 76.595 114.940 ;
        RECT 102.185 114.415 102.355 114.940 ;
        RECT 127.945 114.415 128.115 114.940 ;
      LAYER nwell ;
        RECT 50.330 111.125 139.490 113.955 ;
      LAYER pwell ;
        RECT 63.545 110.140 63.715 110.665 ;
        RECT 89.305 110.140 89.475 110.665 ;
        RECT 115.065 110.140 115.235 110.665 ;
        RECT 50.665 109.735 50.835 109.905 ;
        RECT 52.045 109.735 52.215 109.905 ;
        RECT 57.565 109.735 57.735 109.905 ;
        RECT 63.085 109.875 63.255 109.905 ;
        RECT 63.080 109.765 63.255 109.875 ;
        RECT 63.085 109.735 63.255 109.765 ;
        RECT 64.005 109.735 64.175 109.905 ;
        RECT 64.920 109.765 65.040 109.875 ;
        RECT 65.385 109.735 65.555 109.905 ;
        RECT 66.765 109.735 66.935 109.905 ;
        RECT 68.605 109.735 68.775 109.905 ;
        RECT 69.525 109.735 69.695 109.905 ;
        RECT 74.125 109.735 74.295 109.905 ;
        RECT 75.045 109.735 75.215 109.905 ;
        RECT 75.960 109.765 76.080 109.875 ;
        RECT 76.885 109.735 77.055 109.905 ;
        RECT 80.565 109.735 80.735 109.905 ;
        RECT 82.405 109.735 82.575 109.905 ;
        RECT 86.085 109.735 86.255 109.905 ;
        RECT 87.925 109.735 88.095 109.905 ;
        RECT 88.840 109.765 88.960 109.875 ;
        RECT 89.765 109.735 89.935 109.905 ;
        RECT 93.445 109.735 93.615 109.905 ;
        RECT 95.285 109.735 95.455 109.905 ;
        RECT 98.965 109.735 99.135 109.905 ;
        RECT 100.805 109.735 100.975 109.905 ;
        RECT 101.720 109.765 101.840 109.875 ;
        RECT 102.645 109.735 102.815 109.905 ;
        RECT 106.325 109.735 106.495 109.905 ;
        RECT 108.165 109.735 108.335 109.905 ;
        RECT 111.845 109.735 112.015 109.905 ;
        RECT 113.685 109.735 113.855 109.905 ;
        RECT 114.600 109.765 114.720 109.875 ;
        RECT 115.525 109.735 115.695 109.905 ;
        RECT 119.205 109.735 119.375 109.905 ;
        RECT 121.045 109.735 121.215 109.905 ;
        RECT 124.725 109.735 124.895 109.905 ;
        RECT 126.565 109.735 126.735 109.905 ;
        RECT 127.480 109.765 127.600 109.875 ;
        RECT 128.405 109.735 128.575 109.905 ;
        RECT 132.085 109.735 132.255 109.905 ;
        RECT 133.925 109.735 134.095 109.905 ;
        RECT 137.600 109.765 137.720 109.875 ;
        RECT 138.985 109.735 139.155 109.905 ;
        RECT 76.425 108.975 76.595 109.500 ;
        RECT 102.185 108.975 102.355 109.500 ;
        RECT 127.945 108.975 128.115 109.500 ;
      LAYER nwell ;
        RECT 50.330 105.685 139.490 108.515 ;
      LAYER pwell ;
        RECT 63.545 104.700 63.715 105.225 ;
        RECT 89.305 104.700 89.475 105.225 ;
        RECT 115.065 104.700 115.235 105.225 ;
        RECT 50.665 104.295 50.835 104.465 ;
        RECT 52.045 104.295 52.225 104.465 ;
        RECT 53.425 104.295 53.595 104.465 ;
        RECT 55.720 104.325 55.840 104.435 ;
        RECT 57.105 104.295 57.275 104.465 ;
        RECT 57.560 104.295 57.730 104.465 ;
        RECT 58.955 104.320 59.115 104.430 ;
        RECT 59.870 104.295 60.040 104.465 ;
        RECT 62.160 104.295 62.340 104.465 ;
        RECT 62.635 104.330 62.795 104.440 ;
        RECT 64.005 104.295 64.175 104.465 ;
        RECT 66.305 104.295 66.475 104.465 ;
        RECT 69.525 104.295 69.695 104.465 ;
        RECT 71.825 104.295 71.995 104.465 ;
        RECT 75.045 104.295 75.215 104.465 ;
        RECT 75.515 104.320 75.675 104.430 ;
        RECT 76.885 104.295 77.055 104.465 ;
        RECT 80.565 104.295 80.735 104.465 ;
        RECT 82.405 104.295 82.575 104.465 ;
        RECT 86.085 104.295 86.255 104.465 ;
        RECT 87.925 104.295 88.095 104.465 ;
        RECT 88.840 104.325 88.960 104.435 ;
        RECT 89.765 104.295 89.935 104.465 ;
        RECT 93.445 104.295 93.615 104.465 ;
        RECT 95.285 104.295 95.455 104.465 ;
        RECT 98.965 104.295 99.135 104.465 ;
        RECT 100.805 104.295 100.975 104.465 ;
        RECT 101.720 104.325 101.840 104.435 ;
        RECT 102.645 104.295 102.815 104.465 ;
        RECT 106.325 104.295 106.495 104.465 ;
        RECT 108.165 104.295 108.335 104.465 ;
        RECT 111.845 104.295 112.015 104.465 ;
        RECT 113.685 104.295 113.855 104.465 ;
        RECT 114.600 104.325 114.720 104.435 ;
        RECT 115.525 104.295 115.695 104.465 ;
        RECT 119.205 104.295 119.375 104.465 ;
        RECT 121.045 104.295 121.215 104.465 ;
        RECT 124.725 104.295 124.895 104.465 ;
        RECT 126.565 104.295 126.735 104.465 ;
        RECT 127.480 104.325 127.600 104.435 ;
        RECT 128.405 104.295 128.575 104.465 ;
        RECT 132.085 104.295 132.255 104.465 ;
        RECT 133.925 104.295 134.095 104.465 ;
        RECT 137.600 104.325 137.720 104.435 ;
        RECT 138.985 104.295 139.155 104.465 ;
        RECT 76.425 103.535 76.595 104.060 ;
        RECT 102.185 103.535 102.355 104.060 ;
        RECT 127.945 103.535 128.115 104.060 ;
      LAYER nwell ;
        RECT 50.330 100.245 139.490 103.075 ;
      LAYER pwell ;
        RECT 63.545 99.260 63.715 99.785 ;
        RECT 89.305 99.260 89.475 99.785 ;
        RECT 115.065 99.260 115.235 99.785 ;
        RECT 50.665 98.855 50.835 99.025 ;
        RECT 52.045 98.855 52.225 99.025 ;
        RECT 53.425 98.855 53.595 99.025 ;
        RECT 57.565 98.855 57.735 99.025 ;
        RECT 58.945 98.855 59.115 99.025 ;
        RECT 60.320 98.885 60.440 98.995 ;
        RECT 60.785 98.855 60.955 99.025 ;
        RECT 62.165 98.855 62.335 99.025 ;
        RECT 62.635 98.890 62.795 99.000 ;
        RECT 64.005 98.855 64.175 99.025 ;
        RECT 67.685 98.855 67.855 99.025 ;
        RECT 69.525 98.855 69.695 99.025 ;
        RECT 73.205 98.855 73.375 99.025 ;
        RECT 75.045 98.855 75.215 99.025 ;
        RECT 75.960 98.885 76.080 98.995 ;
        RECT 76.885 98.855 77.055 99.025 ;
        RECT 80.565 98.855 80.735 99.025 ;
        RECT 82.405 98.855 82.575 99.025 ;
        RECT 86.085 98.855 86.255 99.025 ;
        RECT 87.925 98.855 88.095 99.025 ;
        RECT 88.840 98.885 88.960 98.995 ;
        RECT 89.765 98.855 89.935 99.025 ;
        RECT 93.445 98.855 93.615 99.025 ;
        RECT 95.285 98.855 95.455 99.025 ;
        RECT 98.965 98.855 99.135 99.025 ;
        RECT 100.805 98.855 100.975 99.025 ;
        RECT 101.720 98.885 101.840 98.995 ;
        RECT 102.645 98.855 102.815 99.025 ;
        RECT 106.325 98.855 106.495 99.025 ;
        RECT 108.165 98.855 108.335 99.025 ;
        RECT 111.845 98.855 112.015 99.025 ;
        RECT 113.685 98.855 113.855 99.025 ;
        RECT 114.600 98.885 114.720 98.995 ;
        RECT 115.525 98.855 115.695 99.025 ;
        RECT 119.205 98.855 119.375 99.025 ;
        RECT 121.045 98.855 121.215 99.025 ;
        RECT 124.725 98.855 124.895 99.025 ;
        RECT 126.565 98.855 126.735 99.025 ;
        RECT 127.480 98.885 127.600 98.995 ;
        RECT 128.405 98.855 128.575 99.025 ;
        RECT 132.085 98.855 132.255 99.025 ;
        RECT 133.925 98.855 134.095 99.025 ;
        RECT 137.600 98.885 137.720 98.995 ;
        RECT 138.985 98.855 139.155 99.025 ;
        RECT 76.425 98.095 76.595 98.620 ;
        RECT 102.185 98.095 102.355 98.620 ;
        RECT 127.945 98.095 128.115 98.620 ;
      LAYER nwell ;
        RECT 50.330 94.805 139.490 97.635 ;
      LAYER pwell ;
        RECT 63.545 93.820 63.715 94.345 ;
        RECT 89.305 93.820 89.475 94.345 ;
        RECT 115.065 93.820 115.235 94.345 ;
        RECT 50.665 93.415 50.835 93.585 ;
        RECT 52.045 93.415 52.215 93.585 ;
        RECT 55.735 93.440 55.895 93.550 ;
        RECT 57.565 93.415 57.735 93.585 ;
        RECT 60.050 93.415 60.220 93.585 ;
        RECT 61.060 93.415 61.230 93.585 ;
        RECT 61.240 93.445 61.360 93.555 ;
        RECT 62.630 93.415 62.800 93.585 ;
        RECT 63.080 93.445 63.200 93.555 ;
        RECT 64.005 93.415 64.175 93.585 ;
        RECT 64.925 93.415 65.095 93.585 ;
        RECT 66.305 93.415 66.475 93.585 ;
        RECT 67.685 93.415 67.855 93.585 ;
        RECT 69.525 93.415 69.695 93.585 ;
        RECT 73.205 93.415 73.375 93.585 ;
        RECT 75.045 93.415 75.215 93.585 ;
        RECT 75.960 93.445 76.080 93.555 ;
        RECT 76.885 93.415 77.055 93.585 ;
        RECT 80.565 93.415 80.735 93.585 ;
        RECT 82.405 93.415 82.575 93.585 ;
        RECT 86.085 93.415 86.255 93.585 ;
        RECT 87.925 93.415 88.095 93.585 ;
        RECT 88.840 93.445 88.960 93.555 ;
        RECT 89.765 93.415 89.935 93.585 ;
        RECT 93.445 93.415 93.615 93.585 ;
        RECT 95.285 93.415 95.455 93.585 ;
        RECT 98.965 93.415 99.135 93.585 ;
        RECT 100.805 93.415 100.975 93.585 ;
        RECT 101.720 93.445 101.840 93.555 ;
        RECT 102.645 93.415 102.815 93.585 ;
        RECT 106.325 93.415 106.495 93.585 ;
        RECT 108.165 93.415 108.335 93.585 ;
        RECT 111.845 93.415 112.015 93.585 ;
        RECT 113.685 93.415 113.855 93.585 ;
        RECT 114.600 93.445 114.720 93.555 ;
        RECT 115.525 93.415 115.695 93.585 ;
        RECT 119.205 93.415 119.375 93.585 ;
        RECT 121.045 93.415 121.215 93.585 ;
        RECT 124.725 93.415 124.895 93.585 ;
        RECT 126.565 93.415 126.735 93.585 ;
        RECT 127.480 93.445 127.600 93.555 ;
        RECT 128.405 93.415 128.575 93.585 ;
        RECT 132.085 93.415 132.255 93.585 ;
        RECT 133.925 93.415 134.095 93.585 ;
        RECT 137.600 93.445 137.720 93.555 ;
        RECT 138.985 93.415 139.155 93.585 ;
        RECT 76.425 92.655 76.595 93.180 ;
        RECT 102.185 92.655 102.355 93.180 ;
        RECT 127.945 92.655 128.115 93.180 ;
      LAYER nwell ;
        RECT 50.330 89.365 139.490 92.195 ;
      LAYER pwell ;
        RECT 63.545 88.380 63.715 88.905 ;
        RECT 89.305 88.380 89.475 88.905 ;
        RECT 115.065 88.380 115.235 88.905 ;
        RECT 50.665 87.975 50.835 88.145 ;
        RECT 52.045 87.975 52.215 88.145 ;
        RECT 57.565 87.975 57.735 88.145 ;
        RECT 60.335 87.975 60.505 88.145 ;
        RECT 61.705 87.975 61.875 88.145 ;
        RECT 63.085 88.115 63.255 88.145 ;
        RECT 63.080 88.005 63.255 88.115 ;
        RECT 63.085 87.975 63.255 88.005 ;
        RECT 64.005 87.975 64.175 88.145 ;
        RECT 68.605 87.975 68.775 88.145 ;
        RECT 69.525 87.975 69.695 88.145 ;
        RECT 74.125 87.975 74.295 88.145 ;
        RECT 75.045 87.975 75.215 88.145 ;
        RECT 75.960 88.005 76.080 88.115 ;
        RECT 76.885 87.975 77.055 88.145 ;
        RECT 80.565 87.975 80.735 88.145 ;
        RECT 82.405 87.975 82.575 88.145 ;
        RECT 86.085 87.975 86.255 88.145 ;
        RECT 87.925 87.975 88.095 88.145 ;
        RECT 88.840 88.005 88.960 88.115 ;
        RECT 89.765 87.975 89.935 88.145 ;
        RECT 93.445 87.975 93.615 88.145 ;
        RECT 95.285 87.975 95.455 88.145 ;
        RECT 98.965 87.975 99.135 88.145 ;
        RECT 100.805 87.975 100.975 88.145 ;
        RECT 101.720 88.005 101.840 88.115 ;
        RECT 102.645 87.975 102.815 88.145 ;
        RECT 106.325 87.975 106.495 88.145 ;
        RECT 108.165 87.975 108.335 88.145 ;
        RECT 111.845 87.975 112.015 88.145 ;
        RECT 113.685 87.975 113.855 88.145 ;
        RECT 114.600 88.005 114.720 88.115 ;
        RECT 115.525 87.975 115.695 88.145 ;
        RECT 119.205 87.975 119.375 88.145 ;
        RECT 121.045 87.975 121.215 88.145 ;
        RECT 124.725 87.975 124.895 88.145 ;
        RECT 126.565 87.975 126.735 88.145 ;
        RECT 127.480 88.005 127.600 88.115 ;
        RECT 128.405 87.975 128.575 88.145 ;
        RECT 132.085 87.975 132.255 88.145 ;
        RECT 133.925 87.975 134.095 88.145 ;
        RECT 137.600 88.005 137.720 88.115 ;
        RECT 138.985 87.975 139.155 88.145 ;
        RECT 76.425 87.215 76.595 87.740 ;
        RECT 102.185 87.215 102.355 87.740 ;
        RECT 127.945 87.215 128.115 87.740 ;
      LAYER nwell ;
        RECT 50.330 83.925 139.490 86.755 ;
      LAYER pwell ;
        RECT 63.545 82.940 63.715 83.465 ;
        RECT 89.305 82.940 89.475 83.465 ;
        RECT 115.065 82.940 115.235 83.465 ;
        RECT 50.665 82.535 50.835 82.705 ;
        RECT 52.045 82.535 52.215 82.705 ;
        RECT 57.565 82.535 57.735 82.705 ;
        RECT 63.085 82.675 63.255 82.705 ;
        RECT 63.080 82.565 63.255 82.675 ;
        RECT 63.085 82.535 63.255 82.565 ;
        RECT 64.005 82.535 64.175 82.705 ;
        RECT 68.605 82.535 68.775 82.705 ;
        RECT 69.525 82.535 69.695 82.705 ;
        RECT 74.125 82.535 74.295 82.705 ;
        RECT 75.045 82.535 75.215 82.705 ;
        RECT 75.960 82.565 76.080 82.675 ;
        RECT 76.885 82.535 77.055 82.705 ;
        RECT 80.565 82.535 80.735 82.705 ;
        RECT 82.405 82.535 82.575 82.705 ;
        RECT 86.085 82.535 86.255 82.705 ;
        RECT 87.925 82.535 88.095 82.705 ;
        RECT 88.840 82.565 88.960 82.675 ;
        RECT 89.765 82.535 89.935 82.705 ;
        RECT 93.445 82.535 93.615 82.705 ;
        RECT 95.285 82.535 95.455 82.705 ;
        RECT 98.965 82.535 99.135 82.705 ;
        RECT 100.805 82.535 100.975 82.705 ;
        RECT 101.720 82.565 101.840 82.675 ;
        RECT 102.645 82.535 102.815 82.705 ;
        RECT 106.325 82.535 106.495 82.705 ;
        RECT 108.165 82.535 108.335 82.705 ;
        RECT 111.845 82.535 112.015 82.705 ;
        RECT 113.685 82.535 113.855 82.705 ;
        RECT 114.600 82.565 114.720 82.675 ;
        RECT 115.525 82.535 115.695 82.705 ;
        RECT 119.205 82.535 119.375 82.705 ;
        RECT 121.045 82.535 121.215 82.705 ;
        RECT 124.725 82.535 124.895 82.705 ;
        RECT 126.565 82.535 126.735 82.705 ;
        RECT 127.480 82.565 127.600 82.675 ;
        RECT 128.405 82.535 128.575 82.705 ;
        RECT 132.085 82.535 132.255 82.705 ;
        RECT 133.925 82.535 134.095 82.705 ;
        RECT 137.600 82.565 137.720 82.675 ;
        RECT 138.985 82.535 139.155 82.705 ;
        RECT 76.425 81.775 76.595 82.300 ;
        RECT 102.185 81.775 102.355 82.300 ;
        RECT 127.945 81.775 128.115 82.300 ;
      LAYER nwell ;
        RECT 50.330 78.485 139.490 81.315 ;
      LAYER pwell ;
        RECT 63.545 77.500 63.715 78.025 ;
        RECT 89.305 77.500 89.475 78.025 ;
        RECT 115.065 77.500 115.235 78.025 ;
        RECT 50.665 77.095 50.835 77.265 ;
        RECT 52.045 77.095 52.215 77.265 ;
        RECT 57.565 77.095 57.735 77.265 ;
        RECT 63.085 77.235 63.255 77.265 ;
        RECT 63.080 77.125 63.255 77.235 ;
        RECT 63.085 77.095 63.255 77.125 ;
        RECT 64.005 77.095 64.175 77.265 ;
        RECT 68.605 77.095 68.775 77.265 ;
        RECT 69.525 77.095 69.695 77.265 ;
        RECT 74.125 77.095 74.295 77.265 ;
        RECT 75.045 77.095 75.215 77.265 ;
        RECT 75.960 77.125 76.080 77.235 ;
        RECT 76.885 77.095 77.055 77.265 ;
        RECT 80.565 77.095 80.735 77.265 ;
        RECT 82.405 77.095 82.575 77.265 ;
        RECT 86.085 77.095 86.255 77.265 ;
        RECT 87.925 77.095 88.095 77.265 ;
        RECT 88.840 77.125 88.960 77.235 ;
        RECT 89.765 77.095 89.935 77.265 ;
        RECT 93.445 77.095 93.615 77.265 ;
        RECT 95.285 77.095 95.455 77.265 ;
        RECT 98.965 77.095 99.135 77.265 ;
        RECT 100.805 77.095 100.975 77.265 ;
        RECT 101.720 77.125 101.840 77.235 ;
        RECT 102.645 77.095 102.815 77.265 ;
        RECT 106.325 77.095 106.495 77.265 ;
        RECT 108.165 77.095 108.335 77.265 ;
        RECT 111.845 77.095 112.015 77.265 ;
        RECT 113.685 77.095 113.855 77.265 ;
        RECT 114.600 77.125 114.720 77.235 ;
        RECT 115.525 77.095 115.695 77.265 ;
        RECT 119.205 77.095 119.375 77.265 ;
        RECT 121.045 77.095 121.215 77.265 ;
        RECT 124.725 77.095 124.895 77.265 ;
        RECT 126.565 77.095 126.735 77.265 ;
        RECT 127.480 77.125 127.600 77.235 ;
        RECT 128.405 77.095 128.575 77.265 ;
        RECT 132.085 77.095 132.255 77.265 ;
        RECT 133.925 77.095 134.095 77.265 ;
        RECT 137.600 77.125 137.720 77.235 ;
        RECT 138.985 77.095 139.155 77.265 ;
        RECT 76.425 76.335 76.595 76.860 ;
        RECT 102.185 76.335 102.355 76.860 ;
        RECT 127.945 76.335 128.115 76.860 ;
      LAYER nwell ;
        RECT 50.330 73.045 139.490 75.875 ;
      LAYER pwell ;
        RECT 63.545 72.060 63.715 72.585 ;
        RECT 89.305 72.060 89.475 72.585 ;
        RECT 115.065 72.060 115.235 72.585 ;
        RECT 50.665 71.655 50.835 71.825 ;
        RECT 52.045 71.655 52.215 71.825 ;
        RECT 57.565 71.655 57.735 71.825 ;
        RECT 63.085 71.795 63.255 71.825 ;
        RECT 63.080 71.685 63.255 71.795 ;
        RECT 63.085 71.655 63.255 71.685 ;
        RECT 64.005 71.655 64.175 71.825 ;
        RECT 68.605 71.655 68.775 71.825 ;
        RECT 69.525 71.655 69.695 71.825 ;
        RECT 74.125 71.655 74.295 71.825 ;
        RECT 75.045 71.655 75.215 71.825 ;
        RECT 75.960 71.685 76.080 71.795 ;
        RECT 76.885 71.655 77.055 71.825 ;
        RECT 80.565 71.655 80.735 71.825 ;
        RECT 82.405 71.655 82.575 71.825 ;
        RECT 86.085 71.655 86.255 71.825 ;
        RECT 87.925 71.655 88.095 71.825 ;
        RECT 88.840 71.685 88.960 71.795 ;
        RECT 89.765 71.655 89.935 71.825 ;
        RECT 93.445 71.655 93.615 71.825 ;
        RECT 95.285 71.655 95.455 71.825 ;
        RECT 98.965 71.655 99.135 71.825 ;
        RECT 100.805 71.655 100.975 71.825 ;
        RECT 101.720 71.685 101.840 71.795 ;
        RECT 102.645 71.655 102.815 71.825 ;
        RECT 106.325 71.655 106.495 71.825 ;
        RECT 108.165 71.655 108.335 71.825 ;
        RECT 111.845 71.655 112.015 71.825 ;
        RECT 113.685 71.655 113.855 71.825 ;
        RECT 114.600 71.685 114.720 71.795 ;
        RECT 115.525 71.655 115.695 71.825 ;
        RECT 119.205 71.655 119.375 71.825 ;
        RECT 121.045 71.655 121.215 71.825 ;
        RECT 124.725 71.655 124.895 71.825 ;
        RECT 126.565 71.655 126.735 71.825 ;
        RECT 127.480 71.685 127.600 71.795 ;
        RECT 128.405 71.655 128.575 71.825 ;
        RECT 132.085 71.655 132.255 71.825 ;
        RECT 133.925 71.655 134.095 71.825 ;
        RECT 137.600 71.685 137.720 71.795 ;
        RECT 138.985 71.655 139.155 71.825 ;
        RECT 76.425 70.895 76.595 71.420 ;
        RECT 102.185 70.895 102.355 71.420 ;
        RECT 127.945 70.895 128.115 71.420 ;
      LAYER nwell ;
        RECT 50.330 67.605 139.490 70.435 ;
      LAYER pwell ;
        RECT 63.545 66.620 63.715 67.145 ;
        RECT 89.305 66.620 89.475 67.145 ;
        RECT 115.065 66.620 115.235 67.145 ;
        RECT 50.665 66.215 50.835 66.385 ;
        RECT 52.045 66.215 52.215 66.385 ;
        RECT 57.565 66.215 57.735 66.385 ;
        RECT 63.085 66.355 63.255 66.385 ;
        RECT 63.080 66.245 63.255 66.355 ;
        RECT 63.085 66.215 63.255 66.245 ;
        RECT 64.005 66.215 64.175 66.385 ;
        RECT 68.605 66.215 68.775 66.385 ;
        RECT 69.525 66.215 69.695 66.385 ;
        RECT 74.125 66.215 74.295 66.385 ;
        RECT 75.045 66.215 75.215 66.385 ;
        RECT 75.960 66.245 76.080 66.355 ;
        RECT 76.885 66.215 77.055 66.385 ;
        RECT 80.565 66.215 80.735 66.385 ;
        RECT 82.405 66.215 82.575 66.385 ;
        RECT 86.085 66.215 86.255 66.385 ;
        RECT 87.925 66.215 88.095 66.385 ;
        RECT 88.840 66.245 88.960 66.355 ;
        RECT 89.765 66.215 89.935 66.385 ;
        RECT 93.445 66.215 93.615 66.385 ;
        RECT 95.285 66.215 95.455 66.385 ;
        RECT 98.965 66.215 99.135 66.385 ;
        RECT 100.805 66.215 100.975 66.385 ;
        RECT 101.720 66.245 101.840 66.355 ;
        RECT 102.645 66.215 102.815 66.385 ;
        RECT 106.325 66.215 106.495 66.385 ;
        RECT 108.165 66.215 108.335 66.385 ;
        RECT 111.845 66.215 112.015 66.385 ;
        RECT 113.685 66.215 113.855 66.385 ;
        RECT 114.600 66.245 114.720 66.355 ;
        RECT 115.525 66.215 115.695 66.385 ;
        RECT 119.205 66.215 119.375 66.385 ;
        RECT 121.045 66.215 121.215 66.385 ;
        RECT 124.725 66.215 124.895 66.385 ;
        RECT 126.565 66.215 126.735 66.385 ;
        RECT 127.480 66.245 127.600 66.355 ;
        RECT 128.405 66.215 128.575 66.385 ;
        RECT 132.085 66.215 132.255 66.385 ;
        RECT 133.925 66.215 134.095 66.385 ;
        RECT 137.600 66.245 137.720 66.355 ;
        RECT 138.985 66.215 139.155 66.385 ;
        RECT 76.425 65.455 76.595 65.980 ;
        RECT 102.185 65.455 102.355 65.980 ;
        RECT 127.945 65.455 128.115 65.980 ;
      LAYER nwell ;
        RECT 50.330 62.165 139.490 64.995 ;
      LAYER pwell ;
        RECT 63.545 61.180 63.715 61.705 ;
        RECT 76.425 61.180 76.595 61.705 ;
        RECT 89.305 61.180 89.475 61.705 ;
        RECT 102.185 61.180 102.355 61.705 ;
        RECT 115.065 61.180 115.235 61.705 ;
        RECT 127.945 61.180 128.115 61.705 ;
        RECT 50.665 60.775 50.835 60.945 ;
        RECT 52.045 60.775 52.215 60.945 ;
        RECT 57.565 60.775 57.735 60.945 ;
        RECT 63.080 60.805 63.200 60.915 ;
        RECT 64.005 60.775 64.175 60.945 ;
        RECT 69.525 60.775 69.695 60.945 ;
        RECT 75.045 60.775 75.215 60.945 ;
        RECT 76.885 60.775 77.055 60.945 ;
        RECT 82.405 60.775 82.575 60.945 ;
        RECT 87.925 60.775 88.095 60.945 ;
        RECT 89.765 60.775 89.935 60.945 ;
        RECT 95.285 60.775 95.455 60.945 ;
        RECT 100.805 60.775 100.975 60.945 ;
        RECT 102.645 60.775 102.815 60.945 ;
        RECT 108.165 60.775 108.335 60.945 ;
        RECT 113.685 60.775 113.855 60.945 ;
        RECT 115.525 60.775 115.695 60.945 ;
        RECT 121.045 60.775 121.215 60.945 ;
        RECT 126.565 60.775 126.735 60.945 ;
        RECT 128.405 60.775 128.575 60.945 ;
        RECT 133.925 60.775 134.095 60.945 ;
        RECT 137.600 60.805 137.720 60.915 ;
        RECT 138.985 60.775 139.155 60.945 ;
      LAYER li1 ;
        RECT 50.520 136.935 139.300 137.105 ;
        RECT 50.605 136.185 51.815 136.935 ;
        RECT 51.985 136.390 57.330 136.935 ;
        RECT 57.505 136.390 62.850 136.935 ;
        RECT 50.605 135.645 51.125 136.185 ;
        RECT 51.295 135.475 51.815 136.015 ;
        RECT 53.570 135.560 53.910 136.390 ;
        RECT 50.605 134.385 51.815 135.475 ;
        RECT 55.390 134.820 55.740 136.070 ;
        RECT 59.090 135.560 59.430 136.390 ;
        RECT 63.485 136.210 63.775 136.935 ;
        RECT 63.945 136.390 69.290 136.935 ;
        RECT 69.465 136.390 74.810 136.935 ;
        RECT 60.910 134.820 61.260 136.070 ;
        RECT 65.530 135.560 65.870 136.390 ;
        RECT 51.985 134.385 57.330 134.820 ;
        RECT 57.505 134.385 62.850 134.820 ;
        RECT 63.485 134.385 63.775 135.550 ;
        RECT 67.350 134.820 67.700 136.070 ;
        RECT 71.050 135.560 71.390 136.390 ;
        RECT 74.985 136.185 76.195 136.935 ;
        RECT 76.365 136.210 76.655 136.935 ;
        RECT 76.825 136.390 82.170 136.935 ;
        RECT 82.345 136.390 87.690 136.935 ;
        RECT 72.870 134.820 73.220 136.070 ;
        RECT 74.985 135.645 75.505 136.185 ;
        RECT 75.675 135.475 76.195 136.015 ;
        RECT 78.410 135.560 78.750 136.390 ;
        RECT 63.945 134.385 69.290 134.820 ;
        RECT 69.465 134.385 74.810 134.820 ;
        RECT 74.985 134.385 76.195 135.475 ;
        RECT 76.365 134.385 76.655 135.550 ;
        RECT 80.230 134.820 80.580 136.070 ;
        RECT 83.930 135.560 84.270 136.390 ;
        RECT 87.865 136.185 89.075 136.935 ;
        RECT 89.245 136.210 89.535 136.935 ;
        RECT 89.705 136.390 95.050 136.935 ;
        RECT 95.225 136.390 100.570 136.935 ;
        RECT 85.750 134.820 86.100 136.070 ;
        RECT 87.865 135.645 88.385 136.185 ;
        RECT 88.555 135.475 89.075 136.015 ;
        RECT 91.290 135.560 91.630 136.390 ;
        RECT 76.825 134.385 82.170 134.820 ;
        RECT 82.345 134.385 87.690 134.820 ;
        RECT 87.865 134.385 89.075 135.475 ;
        RECT 89.245 134.385 89.535 135.550 ;
        RECT 93.110 134.820 93.460 136.070 ;
        RECT 96.810 135.560 97.150 136.390 ;
        RECT 100.745 136.185 101.955 136.935 ;
        RECT 102.125 136.210 102.415 136.935 ;
        RECT 102.585 136.390 107.930 136.935 ;
        RECT 108.105 136.390 113.450 136.935 ;
        RECT 98.630 134.820 98.980 136.070 ;
        RECT 100.745 135.645 101.265 136.185 ;
        RECT 101.435 135.475 101.955 136.015 ;
        RECT 104.170 135.560 104.510 136.390 ;
        RECT 89.705 134.385 95.050 134.820 ;
        RECT 95.225 134.385 100.570 134.820 ;
        RECT 100.745 134.385 101.955 135.475 ;
        RECT 102.125 134.385 102.415 135.550 ;
        RECT 105.990 134.820 106.340 136.070 ;
        RECT 109.690 135.560 110.030 136.390 ;
        RECT 113.625 136.185 114.835 136.935 ;
        RECT 115.005 136.210 115.295 136.935 ;
        RECT 115.465 136.390 120.810 136.935 ;
        RECT 120.985 136.390 126.330 136.935 ;
        RECT 111.510 134.820 111.860 136.070 ;
        RECT 113.625 135.645 114.145 136.185 ;
        RECT 114.315 135.475 114.835 136.015 ;
        RECT 117.050 135.560 117.390 136.390 ;
        RECT 102.585 134.385 107.930 134.820 ;
        RECT 108.105 134.385 113.450 134.820 ;
        RECT 113.625 134.385 114.835 135.475 ;
        RECT 115.005 134.385 115.295 135.550 ;
        RECT 118.870 134.820 119.220 136.070 ;
        RECT 122.570 135.560 122.910 136.390 ;
        RECT 126.505 136.185 127.715 136.935 ;
        RECT 127.885 136.210 128.175 136.935 ;
        RECT 128.345 136.390 133.690 136.935 ;
        RECT 124.390 134.820 124.740 136.070 ;
        RECT 126.505 135.645 127.025 136.185 ;
        RECT 127.195 135.475 127.715 136.015 ;
        RECT 129.930 135.560 130.270 136.390 ;
        RECT 133.865 136.165 137.375 136.935 ;
        RECT 138.005 136.185 139.215 136.935 ;
        RECT 115.465 134.385 120.810 134.820 ;
        RECT 120.985 134.385 126.330 134.820 ;
        RECT 126.505 134.385 127.715 135.475 ;
        RECT 127.885 134.385 128.175 135.550 ;
        RECT 131.750 134.820 132.100 136.070 ;
        RECT 133.865 135.645 135.515 136.165 ;
        RECT 135.685 135.475 137.375 135.995 ;
        RECT 128.345 134.385 133.690 134.820 ;
        RECT 133.865 134.385 137.375 135.475 ;
        RECT 138.005 135.475 138.525 136.015 ;
        RECT 138.695 135.645 139.215 136.185 ;
        RECT 138.005 134.385 139.215 135.475 ;
        RECT 50.520 134.215 139.300 134.385 ;
        RECT 50.605 133.125 51.815 134.215 ;
        RECT 51.985 133.780 57.330 134.215 ;
        RECT 57.505 133.780 62.850 134.215 ;
        RECT 50.605 132.415 51.125 132.955 ;
        RECT 51.295 132.585 51.815 133.125 ;
        RECT 50.605 131.665 51.815 132.415 ;
        RECT 53.570 132.210 53.910 133.040 ;
        RECT 55.390 132.530 55.740 133.780 ;
        RECT 59.090 132.210 59.430 133.040 ;
        RECT 60.910 132.530 61.260 133.780 ;
        RECT 63.485 133.050 63.775 134.215 ;
        RECT 63.945 133.780 69.290 134.215 ;
        RECT 69.465 133.780 74.810 134.215 ;
        RECT 74.985 133.780 80.330 134.215 ;
        RECT 80.505 133.780 85.850 134.215 ;
        RECT 51.985 131.665 57.330 132.210 ;
        RECT 57.505 131.665 62.850 132.210 ;
        RECT 63.485 131.665 63.775 132.390 ;
        RECT 65.530 132.210 65.870 133.040 ;
        RECT 67.350 132.530 67.700 133.780 ;
        RECT 71.050 132.210 71.390 133.040 ;
        RECT 72.870 132.530 73.220 133.780 ;
        RECT 76.570 132.210 76.910 133.040 ;
        RECT 78.390 132.530 78.740 133.780 ;
        RECT 82.090 132.210 82.430 133.040 ;
        RECT 83.910 132.530 84.260 133.780 ;
        RECT 86.025 133.125 88.615 134.215 ;
        RECT 86.025 132.435 87.235 132.955 ;
        RECT 87.405 132.605 88.615 133.125 ;
        RECT 89.245 133.050 89.535 134.215 ;
        RECT 89.705 133.780 95.050 134.215 ;
        RECT 95.225 133.780 100.570 134.215 ;
        RECT 100.745 133.780 106.090 134.215 ;
        RECT 106.265 133.780 111.610 134.215 ;
        RECT 63.945 131.665 69.290 132.210 ;
        RECT 69.465 131.665 74.810 132.210 ;
        RECT 74.985 131.665 80.330 132.210 ;
        RECT 80.505 131.665 85.850 132.210 ;
        RECT 86.025 131.665 88.615 132.435 ;
        RECT 89.245 131.665 89.535 132.390 ;
        RECT 91.290 132.210 91.630 133.040 ;
        RECT 93.110 132.530 93.460 133.780 ;
        RECT 96.810 132.210 97.150 133.040 ;
        RECT 98.630 132.530 98.980 133.780 ;
        RECT 102.330 132.210 102.670 133.040 ;
        RECT 104.150 132.530 104.500 133.780 ;
        RECT 107.850 132.210 108.190 133.040 ;
        RECT 109.670 132.530 110.020 133.780 ;
        RECT 111.785 133.125 114.375 134.215 ;
        RECT 111.785 132.435 112.995 132.955 ;
        RECT 113.165 132.605 114.375 133.125 ;
        RECT 115.005 133.050 115.295 134.215 ;
        RECT 115.465 133.780 120.810 134.215 ;
        RECT 120.985 133.780 126.330 134.215 ;
        RECT 126.505 133.780 131.850 134.215 ;
        RECT 132.025 133.780 137.370 134.215 ;
        RECT 89.705 131.665 95.050 132.210 ;
        RECT 95.225 131.665 100.570 132.210 ;
        RECT 100.745 131.665 106.090 132.210 ;
        RECT 106.265 131.665 111.610 132.210 ;
        RECT 111.785 131.665 114.375 132.435 ;
        RECT 115.005 131.665 115.295 132.390 ;
        RECT 117.050 132.210 117.390 133.040 ;
        RECT 118.870 132.530 119.220 133.780 ;
        RECT 122.570 132.210 122.910 133.040 ;
        RECT 124.390 132.530 124.740 133.780 ;
        RECT 128.090 132.210 128.430 133.040 ;
        RECT 129.910 132.530 130.260 133.780 ;
        RECT 133.610 132.210 133.950 133.040 ;
        RECT 135.430 132.530 135.780 133.780 ;
        RECT 138.005 133.125 139.215 134.215 ;
        RECT 138.005 132.585 138.525 133.125 ;
        RECT 138.695 132.415 139.215 132.955 ;
        RECT 115.465 131.665 120.810 132.210 ;
        RECT 120.985 131.665 126.330 132.210 ;
        RECT 126.505 131.665 131.850 132.210 ;
        RECT 132.025 131.665 137.370 132.210 ;
        RECT 138.005 131.665 139.215 132.415 ;
        RECT 50.520 131.495 139.300 131.665 ;
        RECT 50.605 130.745 51.815 131.495 ;
        RECT 51.985 130.950 57.330 131.495 ;
        RECT 57.505 130.950 62.850 131.495 ;
        RECT 63.025 130.950 68.370 131.495 ;
        RECT 68.545 130.950 73.890 131.495 ;
        RECT 50.605 130.205 51.125 130.745 ;
        RECT 51.295 130.035 51.815 130.575 ;
        RECT 53.570 130.120 53.910 130.950 ;
        RECT 50.605 128.945 51.815 130.035 ;
        RECT 55.390 129.380 55.740 130.630 ;
        RECT 59.090 130.120 59.430 130.950 ;
        RECT 60.910 129.380 61.260 130.630 ;
        RECT 64.610 130.120 64.950 130.950 ;
        RECT 66.430 129.380 66.780 130.630 ;
        RECT 70.130 130.120 70.470 130.950 ;
        RECT 74.065 130.725 75.735 131.495 ;
        RECT 76.365 130.770 76.655 131.495 ;
        RECT 76.825 130.950 82.170 131.495 ;
        RECT 82.345 130.950 87.690 131.495 ;
        RECT 87.865 130.950 93.210 131.495 ;
        RECT 93.385 130.950 98.730 131.495 ;
        RECT 71.950 129.380 72.300 130.630 ;
        RECT 74.065 130.205 74.815 130.725 ;
        RECT 74.985 130.035 75.735 130.555 ;
        RECT 78.410 130.120 78.750 130.950 ;
        RECT 51.985 128.945 57.330 129.380 ;
        RECT 57.505 128.945 62.850 129.380 ;
        RECT 63.025 128.945 68.370 129.380 ;
        RECT 68.545 128.945 73.890 129.380 ;
        RECT 74.065 128.945 75.735 130.035 ;
        RECT 76.365 128.945 76.655 130.110 ;
        RECT 80.230 129.380 80.580 130.630 ;
        RECT 83.930 130.120 84.270 130.950 ;
        RECT 85.750 129.380 86.100 130.630 ;
        RECT 89.450 130.120 89.790 130.950 ;
        RECT 91.270 129.380 91.620 130.630 ;
        RECT 94.970 130.120 95.310 130.950 ;
        RECT 98.905 130.725 101.495 131.495 ;
        RECT 102.125 130.770 102.415 131.495 ;
        RECT 102.585 130.950 107.930 131.495 ;
        RECT 108.105 130.950 113.450 131.495 ;
        RECT 113.625 130.950 118.970 131.495 ;
        RECT 119.145 130.950 124.490 131.495 ;
        RECT 96.790 129.380 97.140 130.630 ;
        RECT 98.905 130.205 100.115 130.725 ;
        RECT 100.285 130.035 101.495 130.555 ;
        RECT 104.170 130.120 104.510 130.950 ;
        RECT 76.825 128.945 82.170 129.380 ;
        RECT 82.345 128.945 87.690 129.380 ;
        RECT 87.865 128.945 93.210 129.380 ;
        RECT 93.385 128.945 98.730 129.380 ;
        RECT 98.905 128.945 101.495 130.035 ;
        RECT 102.125 128.945 102.415 130.110 ;
        RECT 105.990 129.380 106.340 130.630 ;
        RECT 109.690 130.120 110.030 130.950 ;
        RECT 111.510 129.380 111.860 130.630 ;
        RECT 115.210 130.120 115.550 130.950 ;
        RECT 117.030 129.380 117.380 130.630 ;
        RECT 120.730 130.120 121.070 130.950 ;
        RECT 124.665 130.725 127.255 131.495 ;
        RECT 127.885 130.770 128.175 131.495 ;
        RECT 128.345 130.950 133.690 131.495 ;
        RECT 122.550 129.380 122.900 130.630 ;
        RECT 124.665 130.205 125.875 130.725 ;
        RECT 126.045 130.035 127.255 130.555 ;
        RECT 129.930 130.120 130.270 130.950 ;
        RECT 133.865 130.725 137.375 131.495 ;
        RECT 138.005 130.745 139.215 131.495 ;
        RECT 102.585 128.945 107.930 129.380 ;
        RECT 108.105 128.945 113.450 129.380 ;
        RECT 113.625 128.945 118.970 129.380 ;
        RECT 119.145 128.945 124.490 129.380 ;
        RECT 124.665 128.945 127.255 130.035 ;
        RECT 127.885 128.945 128.175 130.110 ;
        RECT 131.750 129.380 132.100 130.630 ;
        RECT 133.865 130.205 135.515 130.725 ;
        RECT 135.685 130.035 137.375 130.555 ;
        RECT 128.345 128.945 133.690 129.380 ;
        RECT 133.865 128.945 137.375 130.035 ;
        RECT 138.005 130.035 138.525 130.575 ;
        RECT 138.695 130.205 139.215 130.745 ;
        RECT 138.005 128.945 139.215 130.035 ;
        RECT 50.520 128.775 139.300 128.945 ;
        RECT 50.605 127.685 51.815 128.775 ;
        RECT 51.985 128.340 57.330 128.775 ;
        RECT 57.505 128.340 62.850 128.775 ;
        RECT 50.605 126.975 51.125 127.515 ;
        RECT 51.295 127.145 51.815 127.685 ;
        RECT 50.605 126.225 51.815 126.975 ;
        RECT 53.570 126.770 53.910 127.600 ;
        RECT 55.390 127.090 55.740 128.340 ;
        RECT 59.090 126.770 59.430 127.600 ;
        RECT 60.910 127.090 61.260 128.340 ;
        RECT 63.485 127.610 63.775 128.775 ;
        RECT 63.945 128.340 69.290 128.775 ;
        RECT 69.465 128.340 74.810 128.775 ;
        RECT 74.985 128.340 80.330 128.775 ;
        RECT 80.505 128.340 85.850 128.775 ;
        RECT 51.985 126.225 57.330 126.770 ;
        RECT 57.505 126.225 62.850 126.770 ;
        RECT 63.485 126.225 63.775 126.950 ;
        RECT 65.530 126.770 65.870 127.600 ;
        RECT 67.350 127.090 67.700 128.340 ;
        RECT 71.050 126.770 71.390 127.600 ;
        RECT 72.870 127.090 73.220 128.340 ;
        RECT 76.570 126.770 76.910 127.600 ;
        RECT 78.390 127.090 78.740 128.340 ;
        RECT 82.090 126.770 82.430 127.600 ;
        RECT 83.910 127.090 84.260 128.340 ;
        RECT 86.025 127.685 88.615 128.775 ;
        RECT 86.025 126.995 87.235 127.515 ;
        RECT 87.405 127.165 88.615 127.685 ;
        RECT 89.245 127.610 89.535 128.775 ;
        RECT 89.705 128.340 95.050 128.775 ;
        RECT 95.225 128.340 100.570 128.775 ;
        RECT 100.745 128.340 106.090 128.775 ;
        RECT 106.265 128.340 111.610 128.775 ;
        RECT 63.945 126.225 69.290 126.770 ;
        RECT 69.465 126.225 74.810 126.770 ;
        RECT 74.985 126.225 80.330 126.770 ;
        RECT 80.505 126.225 85.850 126.770 ;
        RECT 86.025 126.225 88.615 126.995 ;
        RECT 89.245 126.225 89.535 126.950 ;
        RECT 91.290 126.770 91.630 127.600 ;
        RECT 93.110 127.090 93.460 128.340 ;
        RECT 96.810 126.770 97.150 127.600 ;
        RECT 98.630 127.090 98.980 128.340 ;
        RECT 102.330 126.770 102.670 127.600 ;
        RECT 104.150 127.090 104.500 128.340 ;
        RECT 107.850 126.770 108.190 127.600 ;
        RECT 109.670 127.090 110.020 128.340 ;
        RECT 111.785 127.685 114.375 128.775 ;
        RECT 111.785 126.995 112.995 127.515 ;
        RECT 113.165 127.165 114.375 127.685 ;
        RECT 115.005 127.610 115.295 128.775 ;
        RECT 115.465 128.340 120.810 128.775 ;
        RECT 120.985 128.340 126.330 128.775 ;
        RECT 126.505 128.340 131.850 128.775 ;
        RECT 132.025 128.340 137.370 128.775 ;
        RECT 89.705 126.225 95.050 126.770 ;
        RECT 95.225 126.225 100.570 126.770 ;
        RECT 100.745 126.225 106.090 126.770 ;
        RECT 106.265 126.225 111.610 126.770 ;
        RECT 111.785 126.225 114.375 126.995 ;
        RECT 115.005 126.225 115.295 126.950 ;
        RECT 117.050 126.770 117.390 127.600 ;
        RECT 118.870 127.090 119.220 128.340 ;
        RECT 122.570 126.770 122.910 127.600 ;
        RECT 124.390 127.090 124.740 128.340 ;
        RECT 128.090 126.770 128.430 127.600 ;
        RECT 129.910 127.090 130.260 128.340 ;
        RECT 133.610 126.770 133.950 127.600 ;
        RECT 135.430 127.090 135.780 128.340 ;
        RECT 138.005 127.685 139.215 128.775 ;
        RECT 138.005 127.145 138.525 127.685 ;
        RECT 138.695 126.975 139.215 127.515 ;
        RECT 115.465 126.225 120.810 126.770 ;
        RECT 120.985 126.225 126.330 126.770 ;
        RECT 126.505 126.225 131.850 126.770 ;
        RECT 132.025 126.225 137.370 126.770 ;
        RECT 138.005 126.225 139.215 126.975 ;
        RECT 50.520 126.055 139.300 126.225 ;
        RECT 50.605 125.305 51.815 126.055 ;
        RECT 51.985 125.510 57.330 126.055 ;
        RECT 57.505 125.510 62.850 126.055 ;
        RECT 63.025 125.510 68.370 126.055 ;
        RECT 68.545 125.510 73.890 126.055 ;
        RECT 50.605 124.765 51.125 125.305 ;
        RECT 51.295 124.595 51.815 125.135 ;
        RECT 53.570 124.680 53.910 125.510 ;
        RECT 50.605 123.505 51.815 124.595 ;
        RECT 55.390 123.940 55.740 125.190 ;
        RECT 59.090 124.680 59.430 125.510 ;
        RECT 60.910 123.940 61.260 125.190 ;
        RECT 64.610 124.680 64.950 125.510 ;
        RECT 66.430 123.940 66.780 125.190 ;
        RECT 70.130 124.680 70.470 125.510 ;
        RECT 74.065 125.285 75.735 126.055 ;
        RECT 76.365 125.330 76.655 126.055 ;
        RECT 76.825 125.510 82.170 126.055 ;
        RECT 82.345 125.510 87.690 126.055 ;
        RECT 87.865 125.510 93.210 126.055 ;
        RECT 93.385 125.510 98.730 126.055 ;
        RECT 71.950 123.940 72.300 125.190 ;
        RECT 74.065 124.765 74.815 125.285 ;
        RECT 74.985 124.595 75.735 125.115 ;
        RECT 78.410 124.680 78.750 125.510 ;
        RECT 51.985 123.505 57.330 123.940 ;
        RECT 57.505 123.505 62.850 123.940 ;
        RECT 63.025 123.505 68.370 123.940 ;
        RECT 68.545 123.505 73.890 123.940 ;
        RECT 74.065 123.505 75.735 124.595 ;
        RECT 76.365 123.505 76.655 124.670 ;
        RECT 80.230 123.940 80.580 125.190 ;
        RECT 83.930 124.680 84.270 125.510 ;
        RECT 85.750 123.940 86.100 125.190 ;
        RECT 89.450 124.680 89.790 125.510 ;
        RECT 91.270 123.940 91.620 125.190 ;
        RECT 94.970 124.680 95.310 125.510 ;
        RECT 98.905 125.285 101.495 126.055 ;
        RECT 102.125 125.330 102.415 126.055 ;
        RECT 102.585 125.510 107.930 126.055 ;
        RECT 108.105 125.510 113.450 126.055 ;
        RECT 113.625 125.510 118.970 126.055 ;
        RECT 119.145 125.510 124.490 126.055 ;
        RECT 96.790 123.940 97.140 125.190 ;
        RECT 98.905 124.765 100.115 125.285 ;
        RECT 100.285 124.595 101.495 125.115 ;
        RECT 104.170 124.680 104.510 125.510 ;
        RECT 76.825 123.505 82.170 123.940 ;
        RECT 82.345 123.505 87.690 123.940 ;
        RECT 87.865 123.505 93.210 123.940 ;
        RECT 93.385 123.505 98.730 123.940 ;
        RECT 98.905 123.505 101.495 124.595 ;
        RECT 102.125 123.505 102.415 124.670 ;
        RECT 105.990 123.940 106.340 125.190 ;
        RECT 109.690 124.680 110.030 125.510 ;
        RECT 111.510 123.940 111.860 125.190 ;
        RECT 115.210 124.680 115.550 125.510 ;
        RECT 117.030 123.940 117.380 125.190 ;
        RECT 120.730 124.680 121.070 125.510 ;
        RECT 124.665 125.285 127.255 126.055 ;
        RECT 127.885 125.330 128.175 126.055 ;
        RECT 128.345 125.510 133.690 126.055 ;
        RECT 122.550 123.940 122.900 125.190 ;
        RECT 124.665 124.765 125.875 125.285 ;
        RECT 126.045 124.595 127.255 125.115 ;
        RECT 129.930 124.680 130.270 125.510 ;
        RECT 133.865 125.285 137.375 126.055 ;
        RECT 138.005 125.305 139.215 126.055 ;
        RECT 102.585 123.505 107.930 123.940 ;
        RECT 108.105 123.505 113.450 123.940 ;
        RECT 113.625 123.505 118.970 123.940 ;
        RECT 119.145 123.505 124.490 123.940 ;
        RECT 124.665 123.505 127.255 124.595 ;
        RECT 127.885 123.505 128.175 124.670 ;
        RECT 131.750 123.940 132.100 125.190 ;
        RECT 133.865 124.765 135.515 125.285 ;
        RECT 135.685 124.595 137.375 125.115 ;
        RECT 128.345 123.505 133.690 123.940 ;
        RECT 133.865 123.505 137.375 124.595 ;
        RECT 138.005 124.595 138.525 125.135 ;
        RECT 138.695 124.765 139.215 125.305 ;
        RECT 138.005 123.505 139.215 124.595 ;
        RECT 50.520 123.335 139.300 123.505 ;
        RECT 50.605 122.245 51.815 123.335 ;
        RECT 51.985 122.900 57.330 123.335 ;
        RECT 57.505 122.900 62.850 123.335 ;
        RECT 50.605 121.535 51.125 122.075 ;
        RECT 51.295 121.705 51.815 122.245 ;
        RECT 50.605 120.785 51.815 121.535 ;
        RECT 53.570 121.330 53.910 122.160 ;
        RECT 55.390 121.650 55.740 122.900 ;
        RECT 59.090 121.330 59.430 122.160 ;
        RECT 60.910 121.650 61.260 122.900 ;
        RECT 63.485 122.170 63.775 123.335 ;
        RECT 63.945 122.900 69.290 123.335 ;
        RECT 69.465 122.900 74.810 123.335 ;
        RECT 74.985 122.900 80.330 123.335 ;
        RECT 80.505 122.900 85.850 123.335 ;
        RECT 51.985 120.785 57.330 121.330 ;
        RECT 57.505 120.785 62.850 121.330 ;
        RECT 63.485 120.785 63.775 121.510 ;
        RECT 65.530 121.330 65.870 122.160 ;
        RECT 67.350 121.650 67.700 122.900 ;
        RECT 71.050 121.330 71.390 122.160 ;
        RECT 72.870 121.650 73.220 122.900 ;
        RECT 76.570 121.330 76.910 122.160 ;
        RECT 78.390 121.650 78.740 122.900 ;
        RECT 82.090 121.330 82.430 122.160 ;
        RECT 83.910 121.650 84.260 122.900 ;
        RECT 86.025 122.245 88.615 123.335 ;
        RECT 86.025 121.555 87.235 122.075 ;
        RECT 87.405 121.725 88.615 122.245 ;
        RECT 89.245 122.170 89.535 123.335 ;
        RECT 89.705 122.900 95.050 123.335 ;
        RECT 95.225 122.900 100.570 123.335 ;
        RECT 100.745 122.900 106.090 123.335 ;
        RECT 106.265 122.900 111.610 123.335 ;
        RECT 63.945 120.785 69.290 121.330 ;
        RECT 69.465 120.785 74.810 121.330 ;
        RECT 74.985 120.785 80.330 121.330 ;
        RECT 80.505 120.785 85.850 121.330 ;
        RECT 86.025 120.785 88.615 121.555 ;
        RECT 89.245 120.785 89.535 121.510 ;
        RECT 91.290 121.330 91.630 122.160 ;
        RECT 93.110 121.650 93.460 122.900 ;
        RECT 96.810 121.330 97.150 122.160 ;
        RECT 98.630 121.650 98.980 122.900 ;
        RECT 102.330 121.330 102.670 122.160 ;
        RECT 104.150 121.650 104.500 122.900 ;
        RECT 107.850 121.330 108.190 122.160 ;
        RECT 109.670 121.650 110.020 122.900 ;
        RECT 111.785 122.245 114.375 123.335 ;
        RECT 111.785 121.555 112.995 122.075 ;
        RECT 113.165 121.725 114.375 122.245 ;
        RECT 115.005 122.170 115.295 123.335 ;
        RECT 115.465 122.900 120.810 123.335 ;
        RECT 120.985 122.900 126.330 123.335 ;
        RECT 126.505 122.900 131.850 123.335 ;
        RECT 132.025 122.900 137.370 123.335 ;
        RECT 89.705 120.785 95.050 121.330 ;
        RECT 95.225 120.785 100.570 121.330 ;
        RECT 100.745 120.785 106.090 121.330 ;
        RECT 106.265 120.785 111.610 121.330 ;
        RECT 111.785 120.785 114.375 121.555 ;
        RECT 115.005 120.785 115.295 121.510 ;
        RECT 117.050 121.330 117.390 122.160 ;
        RECT 118.870 121.650 119.220 122.900 ;
        RECT 122.570 121.330 122.910 122.160 ;
        RECT 124.390 121.650 124.740 122.900 ;
        RECT 128.090 121.330 128.430 122.160 ;
        RECT 129.910 121.650 130.260 122.900 ;
        RECT 133.610 121.330 133.950 122.160 ;
        RECT 135.430 121.650 135.780 122.900 ;
        RECT 138.005 122.245 139.215 123.335 ;
        RECT 138.005 121.705 138.525 122.245 ;
        RECT 138.695 121.535 139.215 122.075 ;
        RECT 115.465 120.785 120.810 121.330 ;
        RECT 120.985 120.785 126.330 121.330 ;
        RECT 126.505 120.785 131.850 121.330 ;
        RECT 132.025 120.785 137.370 121.330 ;
        RECT 138.005 120.785 139.215 121.535 ;
        RECT 50.520 120.615 139.300 120.785 ;
        RECT 50.605 119.865 51.815 120.615 ;
        RECT 51.985 120.070 57.330 120.615 ;
        RECT 57.505 120.070 62.850 120.615 ;
        RECT 63.025 120.070 68.370 120.615 ;
        RECT 68.545 120.070 73.890 120.615 ;
        RECT 50.605 119.325 51.125 119.865 ;
        RECT 51.295 119.155 51.815 119.695 ;
        RECT 53.570 119.240 53.910 120.070 ;
        RECT 50.605 118.065 51.815 119.155 ;
        RECT 55.390 118.500 55.740 119.750 ;
        RECT 59.090 119.240 59.430 120.070 ;
        RECT 60.910 118.500 61.260 119.750 ;
        RECT 64.610 119.240 64.950 120.070 ;
        RECT 66.430 118.500 66.780 119.750 ;
        RECT 70.130 119.240 70.470 120.070 ;
        RECT 74.065 119.845 75.735 120.615 ;
        RECT 76.365 119.890 76.655 120.615 ;
        RECT 76.825 120.070 82.170 120.615 ;
        RECT 82.345 120.070 87.690 120.615 ;
        RECT 87.865 120.070 93.210 120.615 ;
        RECT 93.385 120.070 98.730 120.615 ;
        RECT 71.950 118.500 72.300 119.750 ;
        RECT 74.065 119.325 74.815 119.845 ;
        RECT 74.985 119.155 75.735 119.675 ;
        RECT 78.410 119.240 78.750 120.070 ;
        RECT 51.985 118.065 57.330 118.500 ;
        RECT 57.505 118.065 62.850 118.500 ;
        RECT 63.025 118.065 68.370 118.500 ;
        RECT 68.545 118.065 73.890 118.500 ;
        RECT 74.065 118.065 75.735 119.155 ;
        RECT 76.365 118.065 76.655 119.230 ;
        RECT 80.230 118.500 80.580 119.750 ;
        RECT 83.930 119.240 84.270 120.070 ;
        RECT 85.750 118.500 86.100 119.750 ;
        RECT 89.450 119.240 89.790 120.070 ;
        RECT 91.270 118.500 91.620 119.750 ;
        RECT 94.970 119.240 95.310 120.070 ;
        RECT 98.905 119.845 101.495 120.615 ;
        RECT 102.125 119.890 102.415 120.615 ;
        RECT 102.585 120.070 107.930 120.615 ;
        RECT 108.105 120.070 113.450 120.615 ;
        RECT 113.625 120.070 118.970 120.615 ;
        RECT 119.145 120.070 124.490 120.615 ;
        RECT 96.790 118.500 97.140 119.750 ;
        RECT 98.905 119.325 100.115 119.845 ;
        RECT 100.285 119.155 101.495 119.675 ;
        RECT 104.170 119.240 104.510 120.070 ;
        RECT 76.825 118.065 82.170 118.500 ;
        RECT 82.345 118.065 87.690 118.500 ;
        RECT 87.865 118.065 93.210 118.500 ;
        RECT 93.385 118.065 98.730 118.500 ;
        RECT 98.905 118.065 101.495 119.155 ;
        RECT 102.125 118.065 102.415 119.230 ;
        RECT 105.990 118.500 106.340 119.750 ;
        RECT 109.690 119.240 110.030 120.070 ;
        RECT 111.510 118.500 111.860 119.750 ;
        RECT 115.210 119.240 115.550 120.070 ;
        RECT 117.030 118.500 117.380 119.750 ;
        RECT 120.730 119.240 121.070 120.070 ;
        RECT 124.665 119.845 127.255 120.615 ;
        RECT 127.885 119.890 128.175 120.615 ;
        RECT 128.345 120.070 133.690 120.615 ;
        RECT 122.550 118.500 122.900 119.750 ;
        RECT 124.665 119.325 125.875 119.845 ;
        RECT 126.045 119.155 127.255 119.675 ;
        RECT 129.930 119.240 130.270 120.070 ;
        RECT 133.865 119.845 137.375 120.615 ;
        RECT 138.005 119.865 139.215 120.615 ;
        RECT 102.585 118.065 107.930 118.500 ;
        RECT 108.105 118.065 113.450 118.500 ;
        RECT 113.625 118.065 118.970 118.500 ;
        RECT 119.145 118.065 124.490 118.500 ;
        RECT 124.665 118.065 127.255 119.155 ;
        RECT 127.885 118.065 128.175 119.230 ;
        RECT 131.750 118.500 132.100 119.750 ;
        RECT 133.865 119.325 135.515 119.845 ;
        RECT 135.685 119.155 137.375 119.675 ;
        RECT 128.345 118.065 133.690 118.500 ;
        RECT 133.865 118.065 137.375 119.155 ;
        RECT 138.005 119.155 138.525 119.695 ;
        RECT 138.695 119.325 139.215 119.865 ;
        RECT 138.005 118.065 139.215 119.155 ;
        RECT 50.520 117.895 139.300 118.065 ;
        RECT 50.605 116.805 51.815 117.895 ;
        RECT 51.985 117.460 57.330 117.895 ;
        RECT 57.505 117.460 62.850 117.895 ;
        RECT 50.605 116.095 51.125 116.635 ;
        RECT 51.295 116.265 51.815 116.805 ;
        RECT 50.605 115.345 51.815 116.095 ;
        RECT 53.570 115.890 53.910 116.720 ;
        RECT 55.390 116.210 55.740 117.460 ;
        RECT 59.090 115.890 59.430 116.720 ;
        RECT 60.910 116.210 61.260 117.460 ;
        RECT 63.485 116.730 63.775 117.895 ;
        RECT 63.945 117.460 69.290 117.895 ;
        RECT 69.465 117.460 74.810 117.895 ;
        RECT 74.985 117.460 80.330 117.895 ;
        RECT 80.505 117.460 85.850 117.895 ;
        RECT 51.985 115.345 57.330 115.890 ;
        RECT 57.505 115.345 62.850 115.890 ;
        RECT 63.485 115.345 63.775 116.070 ;
        RECT 65.530 115.890 65.870 116.720 ;
        RECT 67.350 116.210 67.700 117.460 ;
        RECT 71.050 115.890 71.390 116.720 ;
        RECT 72.870 116.210 73.220 117.460 ;
        RECT 76.570 115.890 76.910 116.720 ;
        RECT 78.390 116.210 78.740 117.460 ;
        RECT 82.090 115.890 82.430 116.720 ;
        RECT 83.910 116.210 84.260 117.460 ;
        RECT 86.025 116.805 88.615 117.895 ;
        RECT 86.025 116.115 87.235 116.635 ;
        RECT 87.405 116.285 88.615 116.805 ;
        RECT 89.245 116.730 89.535 117.895 ;
        RECT 89.705 117.460 95.050 117.895 ;
        RECT 95.225 117.460 100.570 117.895 ;
        RECT 100.745 117.460 106.090 117.895 ;
        RECT 106.265 117.460 111.610 117.895 ;
        RECT 63.945 115.345 69.290 115.890 ;
        RECT 69.465 115.345 74.810 115.890 ;
        RECT 74.985 115.345 80.330 115.890 ;
        RECT 80.505 115.345 85.850 115.890 ;
        RECT 86.025 115.345 88.615 116.115 ;
        RECT 89.245 115.345 89.535 116.070 ;
        RECT 91.290 115.890 91.630 116.720 ;
        RECT 93.110 116.210 93.460 117.460 ;
        RECT 96.810 115.890 97.150 116.720 ;
        RECT 98.630 116.210 98.980 117.460 ;
        RECT 102.330 115.890 102.670 116.720 ;
        RECT 104.150 116.210 104.500 117.460 ;
        RECT 107.850 115.890 108.190 116.720 ;
        RECT 109.670 116.210 110.020 117.460 ;
        RECT 111.785 116.805 114.375 117.895 ;
        RECT 111.785 116.115 112.995 116.635 ;
        RECT 113.165 116.285 114.375 116.805 ;
        RECT 115.005 116.730 115.295 117.895 ;
        RECT 115.465 117.460 120.810 117.895 ;
        RECT 120.985 117.460 126.330 117.895 ;
        RECT 126.505 117.460 131.850 117.895 ;
        RECT 132.025 117.460 137.370 117.895 ;
        RECT 89.705 115.345 95.050 115.890 ;
        RECT 95.225 115.345 100.570 115.890 ;
        RECT 100.745 115.345 106.090 115.890 ;
        RECT 106.265 115.345 111.610 115.890 ;
        RECT 111.785 115.345 114.375 116.115 ;
        RECT 115.005 115.345 115.295 116.070 ;
        RECT 117.050 115.890 117.390 116.720 ;
        RECT 118.870 116.210 119.220 117.460 ;
        RECT 122.570 115.890 122.910 116.720 ;
        RECT 124.390 116.210 124.740 117.460 ;
        RECT 128.090 115.890 128.430 116.720 ;
        RECT 129.910 116.210 130.260 117.460 ;
        RECT 133.610 115.890 133.950 116.720 ;
        RECT 135.430 116.210 135.780 117.460 ;
        RECT 138.005 116.805 139.215 117.895 ;
        RECT 138.005 116.265 138.525 116.805 ;
        RECT 138.695 116.095 139.215 116.635 ;
        RECT 115.465 115.345 120.810 115.890 ;
        RECT 120.985 115.345 126.330 115.890 ;
        RECT 126.505 115.345 131.850 115.890 ;
        RECT 132.025 115.345 137.370 115.890 ;
        RECT 138.005 115.345 139.215 116.095 ;
        RECT 50.520 115.175 139.300 115.345 ;
        RECT 50.605 114.425 51.815 115.175 ;
        RECT 51.985 114.630 57.330 115.175 ;
        RECT 57.505 114.630 62.850 115.175 ;
        RECT 63.025 114.630 68.370 115.175 ;
        RECT 68.545 114.630 73.890 115.175 ;
        RECT 50.605 113.885 51.125 114.425 ;
        RECT 51.295 113.715 51.815 114.255 ;
        RECT 53.570 113.800 53.910 114.630 ;
        RECT 50.605 112.625 51.815 113.715 ;
        RECT 55.390 113.060 55.740 114.310 ;
        RECT 59.090 113.800 59.430 114.630 ;
        RECT 60.910 113.060 61.260 114.310 ;
        RECT 64.610 113.800 64.950 114.630 ;
        RECT 66.430 113.060 66.780 114.310 ;
        RECT 70.130 113.800 70.470 114.630 ;
        RECT 74.065 114.405 75.735 115.175 ;
        RECT 76.365 114.450 76.655 115.175 ;
        RECT 76.825 114.630 82.170 115.175 ;
        RECT 82.345 114.630 87.690 115.175 ;
        RECT 87.865 114.630 93.210 115.175 ;
        RECT 93.385 114.630 98.730 115.175 ;
        RECT 71.950 113.060 72.300 114.310 ;
        RECT 74.065 113.885 74.815 114.405 ;
        RECT 74.985 113.715 75.735 114.235 ;
        RECT 78.410 113.800 78.750 114.630 ;
        RECT 51.985 112.625 57.330 113.060 ;
        RECT 57.505 112.625 62.850 113.060 ;
        RECT 63.025 112.625 68.370 113.060 ;
        RECT 68.545 112.625 73.890 113.060 ;
        RECT 74.065 112.625 75.735 113.715 ;
        RECT 76.365 112.625 76.655 113.790 ;
        RECT 80.230 113.060 80.580 114.310 ;
        RECT 83.930 113.800 84.270 114.630 ;
        RECT 85.750 113.060 86.100 114.310 ;
        RECT 89.450 113.800 89.790 114.630 ;
        RECT 91.270 113.060 91.620 114.310 ;
        RECT 94.970 113.800 95.310 114.630 ;
        RECT 98.905 114.405 101.495 115.175 ;
        RECT 102.125 114.450 102.415 115.175 ;
        RECT 102.585 114.630 107.930 115.175 ;
        RECT 108.105 114.630 113.450 115.175 ;
        RECT 113.625 114.630 118.970 115.175 ;
        RECT 119.145 114.630 124.490 115.175 ;
        RECT 96.790 113.060 97.140 114.310 ;
        RECT 98.905 113.885 100.115 114.405 ;
        RECT 100.285 113.715 101.495 114.235 ;
        RECT 104.170 113.800 104.510 114.630 ;
        RECT 76.825 112.625 82.170 113.060 ;
        RECT 82.345 112.625 87.690 113.060 ;
        RECT 87.865 112.625 93.210 113.060 ;
        RECT 93.385 112.625 98.730 113.060 ;
        RECT 98.905 112.625 101.495 113.715 ;
        RECT 102.125 112.625 102.415 113.790 ;
        RECT 105.990 113.060 106.340 114.310 ;
        RECT 109.690 113.800 110.030 114.630 ;
        RECT 111.510 113.060 111.860 114.310 ;
        RECT 115.210 113.800 115.550 114.630 ;
        RECT 117.030 113.060 117.380 114.310 ;
        RECT 120.730 113.800 121.070 114.630 ;
        RECT 124.665 114.405 127.255 115.175 ;
        RECT 127.885 114.450 128.175 115.175 ;
        RECT 128.345 114.630 133.690 115.175 ;
        RECT 122.550 113.060 122.900 114.310 ;
        RECT 124.665 113.885 125.875 114.405 ;
        RECT 126.045 113.715 127.255 114.235 ;
        RECT 129.930 113.800 130.270 114.630 ;
        RECT 133.865 114.405 137.375 115.175 ;
        RECT 138.005 114.425 139.215 115.175 ;
        RECT 102.585 112.625 107.930 113.060 ;
        RECT 108.105 112.625 113.450 113.060 ;
        RECT 113.625 112.625 118.970 113.060 ;
        RECT 119.145 112.625 124.490 113.060 ;
        RECT 124.665 112.625 127.255 113.715 ;
        RECT 127.885 112.625 128.175 113.790 ;
        RECT 131.750 113.060 132.100 114.310 ;
        RECT 133.865 113.885 135.515 114.405 ;
        RECT 135.685 113.715 137.375 114.235 ;
        RECT 128.345 112.625 133.690 113.060 ;
        RECT 133.865 112.625 137.375 113.715 ;
        RECT 138.005 113.715 138.525 114.255 ;
        RECT 138.695 113.885 139.215 114.425 ;
        RECT 138.005 112.625 139.215 113.715 ;
        RECT 50.520 112.455 139.300 112.625 ;
        RECT 50.605 111.365 51.815 112.455 ;
        RECT 51.985 112.020 57.330 112.455 ;
        RECT 57.505 112.020 62.850 112.455 ;
        RECT 50.605 110.655 51.125 111.195 ;
        RECT 51.295 110.825 51.815 111.365 ;
        RECT 50.605 109.905 51.815 110.655 ;
        RECT 53.570 110.450 53.910 111.280 ;
        RECT 55.390 110.770 55.740 112.020 ;
        RECT 59.090 110.450 59.430 111.280 ;
        RECT 60.910 110.770 61.260 112.020 ;
        RECT 63.485 111.290 63.775 112.455 ;
        RECT 63.945 112.020 69.290 112.455 ;
        RECT 69.465 112.020 74.810 112.455 ;
        RECT 74.985 112.020 80.330 112.455 ;
        RECT 80.505 112.020 85.850 112.455 ;
        RECT 51.985 109.905 57.330 110.450 ;
        RECT 57.505 109.905 62.850 110.450 ;
        RECT 63.485 109.905 63.775 110.630 ;
        RECT 65.530 110.450 65.870 111.280 ;
        RECT 67.350 110.770 67.700 112.020 ;
        RECT 71.050 110.450 71.390 111.280 ;
        RECT 72.870 110.770 73.220 112.020 ;
        RECT 76.570 110.450 76.910 111.280 ;
        RECT 78.390 110.770 78.740 112.020 ;
        RECT 82.090 110.450 82.430 111.280 ;
        RECT 83.910 110.770 84.260 112.020 ;
        RECT 86.025 111.365 88.615 112.455 ;
        RECT 86.025 110.675 87.235 111.195 ;
        RECT 87.405 110.845 88.615 111.365 ;
        RECT 89.245 111.290 89.535 112.455 ;
        RECT 89.705 112.020 95.050 112.455 ;
        RECT 95.225 112.020 100.570 112.455 ;
        RECT 100.745 112.020 106.090 112.455 ;
        RECT 106.265 112.020 111.610 112.455 ;
        RECT 63.945 109.905 69.290 110.450 ;
        RECT 69.465 109.905 74.810 110.450 ;
        RECT 74.985 109.905 80.330 110.450 ;
        RECT 80.505 109.905 85.850 110.450 ;
        RECT 86.025 109.905 88.615 110.675 ;
        RECT 89.245 109.905 89.535 110.630 ;
        RECT 91.290 110.450 91.630 111.280 ;
        RECT 93.110 110.770 93.460 112.020 ;
        RECT 96.810 110.450 97.150 111.280 ;
        RECT 98.630 110.770 98.980 112.020 ;
        RECT 102.330 110.450 102.670 111.280 ;
        RECT 104.150 110.770 104.500 112.020 ;
        RECT 107.850 110.450 108.190 111.280 ;
        RECT 109.670 110.770 110.020 112.020 ;
        RECT 111.785 111.365 114.375 112.455 ;
        RECT 111.785 110.675 112.995 111.195 ;
        RECT 113.165 110.845 114.375 111.365 ;
        RECT 115.005 111.290 115.295 112.455 ;
        RECT 115.465 112.020 120.810 112.455 ;
        RECT 120.985 112.020 126.330 112.455 ;
        RECT 126.505 112.020 131.850 112.455 ;
        RECT 132.025 112.020 137.370 112.455 ;
        RECT 89.705 109.905 95.050 110.450 ;
        RECT 95.225 109.905 100.570 110.450 ;
        RECT 100.745 109.905 106.090 110.450 ;
        RECT 106.265 109.905 111.610 110.450 ;
        RECT 111.785 109.905 114.375 110.675 ;
        RECT 115.005 109.905 115.295 110.630 ;
        RECT 117.050 110.450 117.390 111.280 ;
        RECT 118.870 110.770 119.220 112.020 ;
        RECT 122.570 110.450 122.910 111.280 ;
        RECT 124.390 110.770 124.740 112.020 ;
        RECT 128.090 110.450 128.430 111.280 ;
        RECT 129.910 110.770 130.260 112.020 ;
        RECT 133.610 110.450 133.950 111.280 ;
        RECT 135.430 110.770 135.780 112.020 ;
        RECT 138.005 111.365 139.215 112.455 ;
        RECT 138.005 110.825 138.525 111.365 ;
        RECT 138.695 110.655 139.215 111.195 ;
        RECT 115.465 109.905 120.810 110.450 ;
        RECT 120.985 109.905 126.330 110.450 ;
        RECT 126.505 109.905 131.850 110.450 ;
        RECT 132.025 109.905 137.370 110.450 ;
        RECT 138.005 109.905 139.215 110.655 ;
        RECT 50.520 109.735 139.300 109.905 ;
        RECT 50.605 108.985 51.815 109.735 ;
        RECT 51.985 109.190 57.330 109.735 ;
        RECT 57.505 109.190 62.850 109.735 ;
        RECT 50.605 108.445 51.125 108.985 ;
        RECT 51.295 108.275 51.815 108.815 ;
        RECT 53.570 108.360 53.910 109.190 ;
        RECT 50.605 107.185 51.815 108.275 ;
        RECT 55.390 107.620 55.740 108.870 ;
        RECT 59.090 108.360 59.430 109.190 ;
        RECT 63.025 108.965 64.695 109.735 ;
        RECT 60.910 107.620 61.260 108.870 ;
        RECT 63.025 108.445 63.775 108.965 ;
        RECT 65.365 108.915 65.595 109.735 ;
        RECT 65.765 108.935 66.095 109.565 ;
        RECT 63.945 108.275 64.695 108.795 ;
        RECT 65.345 108.495 65.675 108.745 ;
        RECT 65.845 108.335 66.095 108.935 ;
        RECT 66.265 108.915 66.475 109.735 ;
        RECT 66.795 109.185 66.965 109.565 ;
        RECT 67.180 109.355 67.510 109.735 ;
        RECT 66.795 109.015 67.510 109.185 ;
        RECT 66.705 108.465 67.060 108.835 ;
        RECT 67.340 108.825 67.510 109.015 ;
        RECT 67.680 108.990 67.935 109.565 ;
        RECT 67.340 108.495 67.595 108.825 ;
        RECT 51.985 107.185 57.330 107.620 ;
        RECT 57.505 107.185 62.850 107.620 ;
        RECT 63.025 107.185 64.695 108.275 ;
        RECT 65.365 107.185 65.595 108.325 ;
        RECT 65.765 107.355 66.095 108.335 ;
        RECT 66.265 107.185 66.475 108.325 ;
        RECT 67.340 108.285 67.510 108.495 ;
        RECT 66.795 108.115 67.510 108.285 ;
        RECT 67.765 108.260 67.935 108.990 ;
        RECT 68.110 108.895 68.370 109.735 ;
        RECT 68.545 109.190 73.890 109.735 ;
        RECT 70.130 108.360 70.470 109.190 ;
        RECT 74.065 108.965 75.735 109.735 ;
        RECT 76.365 109.010 76.655 109.735 ;
        RECT 76.825 109.190 82.170 109.735 ;
        RECT 82.345 109.190 87.690 109.735 ;
        RECT 87.865 109.190 93.210 109.735 ;
        RECT 93.385 109.190 98.730 109.735 ;
        RECT 66.795 107.355 66.965 108.115 ;
        RECT 67.180 107.185 67.510 107.945 ;
        RECT 67.680 107.355 67.935 108.260 ;
        RECT 68.110 107.185 68.370 108.335 ;
        RECT 71.950 107.620 72.300 108.870 ;
        RECT 74.065 108.445 74.815 108.965 ;
        RECT 74.985 108.275 75.735 108.795 ;
        RECT 78.410 108.360 78.750 109.190 ;
        RECT 68.545 107.185 73.890 107.620 ;
        RECT 74.065 107.185 75.735 108.275 ;
        RECT 76.365 107.185 76.655 108.350 ;
        RECT 80.230 107.620 80.580 108.870 ;
        RECT 83.930 108.360 84.270 109.190 ;
        RECT 85.750 107.620 86.100 108.870 ;
        RECT 89.450 108.360 89.790 109.190 ;
        RECT 91.270 107.620 91.620 108.870 ;
        RECT 94.970 108.360 95.310 109.190 ;
        RECT 98.905 108.965 101.495 109.735 ;
        RECT 102.125 109.010 102.415 109.735 ;
        RECT 102.585 109.190 107.930 109.735 ;
        RECT 108.105 109.190 113.450 109.735 ;
        RECT 113.625 109.190 118.970 109.735 ;
        RECT 119.145 109.190 124.490 109.735 ;
        RECT 96.790 107.620 97.140 108.870 ;
        RECT 98.905 108.445 100.115 108.965 ;
        RECT 100.285 108.275 101.495 108.795 ;
        RECT 104.170 108.360 104.510 109.190 ;
        RECT 76.825 107.185 82.170 107.620 ;
        RECT 82.345 107.185 87.690 107.620 ;
        RECT 87.865 107.185 93.210 107.620 ;
        RECT 93.385 107.185 98.730 107.620 ;
        RECT 98.905 107.185 101.495 108.275 ;
        RECT 102.125 107.185 102.415 108.350 ;
        RECT 105.990 107.620 106.340 108.870 ;
        RECT 109.690 108.360 110.030 109.190 ;
        RECT 111.510 107.620 111.860 108.870 ;
        RECT 115.210 108.360 115.550 109.190 ;
        RECT 117.030 107.620 117.380 108.870 ;
        RECT 120.730 108.360 121.070 109.190 ;
        RECT 124.665 108.965 127.255 109.735 ;
        RECT 127.885 109.010 128.175 109.735 ;
        RECT 128.345 109.190 133.690 109.735 ;
        RECT 122.550 107.620 122.900 108.870 ;
        RECT 124.665 108.445 125.875 108.965 ;
        RECT 126.045 108.275 127.255 108.795 ;
        RECT 129.930 108.360 130.270 109.190 ;
        RECT 133.865 108.965 137.375 109.735 ;
        RECT 138.005 108.985 139.215 109.735 ;
        RECT 102.585 107.185 107.930 107.620 ;
        RECT 108.105 107.185 113.450 107.620 ;
        RECT 113.625 107.185 118.970 107.620 ;
        RECT 119.145 107.185 124.490 107.620 ;
        RECT 124.665 107.185 127.255 108.275 ;
        RECT 127.885 107.185 128.175 108.350 ;
        RECT 131.750 107.620 132.100 108.870 ;
        RECT 133.865 108.445 135.515 108.965 ;
        RECT 135.685 108.275 137.375 108.795 ;
        RECT 128.345 107.185 133.690 107.620 ;
        RECT 133.865 107.185 137.375 108.275 ;
        RECT 138.005 108.275 138.525 108.815 ;
        RECT 138.695 108.445 139.215 108.985 ;
        RECT 138.005 107.185 139.215 108.275 ;
        RECT 50.520 107.015 139.300 107.185 ;
        RECT 50.605 105.925 51.815 107.015 ;
        RECT 51.985 105.925 55.495 107.015 ;
        RECT 50.605 105.215 51.125 105.755 ;
        RECT 51.295 105.385 51.815 105.925 ;
        RECT 51.985 105.235 53.635 105.755 ;
        RECT 53.805 105.405 55.495 105.925 ;
        RECT 56.185 105.875 56.395 107.015 ;
        RECT 56.565 105.865 56.895 106.845 ;
        RECT 57.065 105.875 57.295 107.015 ;
        RECT 57.505 105.875 57.785 107.015 ;
        RECT 57.955 105.865 58.285 106.845 ;
        RECT 58.455 105.875 58.715 107.015 ;
        RECT 58.885 105.875 60.505 106.845 ;
        RECT 60.675 106.555 61.040 107.015 ;
        RECT 61.210 106.385 61.465 106.840 ;
        RECT 61.635 106.555 61.965 107.015 ;
        RECT 62.135 106.385 62.395 106.845 ;
        RECT 60.675 106.180 61.465 106.385 ;
        RECT 50.605 104.465 51.815 105.215 ;
        RECT 51.985 104.465 55.495 105.235 ;
        RECT 56.185 104.465 56.395 105.285 ;
        RECT 56.565 105.265 56.815 105.865 ;
        RECT 58.020 105.825 58.195 105.865 ;
        RECT 56.985 105.455 57.315 105.705 ;
        RECT 57.515 105.435 57.850 105.705 ;
        RECT 56.565 104.635 56.895 105.265 ;
        RECT 57.065 104.465 57.295 105.285 ;
        RECT 58.020 105.265 58.190 105.825 ;
        RECT 58.360 105.455 58.695 105.705 ;
        RECT 57.505 104.465 57.815 105.265 ;
        RECT 58.020 104.635 58.715 105.265 ;
        RECT 58.885 105.205 59.225 105.875 ;
        RECT 60.675 105.705 61.070 106.180 ;
        RECT 61.740 106.165 62.395 106.385 ;
        RECT 59.395 105.375 59.775 105.705 ;
        RECT 59.945 105.455 61.070 105.705 ;
        RECT 61.240 105.455 61.570 106.010 ;
        RECT 59.525 105.285 59.775 105.375 ;
        RECT 58.885 104.635 59.355 105.205 ;
        RECT 59.525 105.115 60.625 105.285 ;
        RECT 59.525 104.465 60.285 104.945 ;
        RECT 60.455 104.845 60.625 105.115 ;
        RECT 60.795 105.265 61.070 105.455 ;
        RECT 60.795 105.015 61.125 105.265 ;
        RECT 61.740 105.205 61.955 106.165 ;
        RECT 62.125 105.375 62.395 105.995 ;
        RECT 63.485 105.850 63.775 107.015 ;
        RECT 63.945 106.580 69.290 107.015 ;
        RECT 69.465 106.580 74.810 107.015 ;
        RECT 74.985 106.580 80.330 107.015 ;
        RECT 80.505 106.580 85.850 107.015 ;
        RECT 61.295 104.995 62.395 105.205 ;
        RECT 61.295 104.845 61.465 104.995 ;
        RECT 60.455 104.635 61.465 104.845 ;
        RECT 61.635 104.465 61.965 104.825 ;
        RECT 62.135 104.660 62.395 104.995 ;
        RECT 63.485 104.465 63.775 105.190 ;
        RECT 65.530 105.010 65.870 105.840 ;
        RECT 67.350 105.330 67.700 106.580 ;
        RECT 71.050 105.010 71.390 105.840 ;
        RECT 72.870 105.330 73.220 106.580 ;
        RECT 76.570 105.010 76.910 105.840 ;
        RECT 78.390 105.330 78.740 106.580 ;
        RECT 82.090 105.010 82.430 105.840 ;
        RECT 83.910 105.330 84.260 106.580 ;
        RECT 86.025 105.925 88.615 107.015 ;
        RECT 86.025 105.235 87.235 105.755 ;
        RECT 87.405 105.405 88.615 105.925 ;
        RECT 89.245 105.850 89.535 107.015 ;
        RECT 89.705 106.580 95.050 107.015 ;
        RECT 95.225 106.580 100.570 107.015 ;
        RECT 100.745 106.580 106.090 107.015 ;
        RECT 106.265 106.580 111.610 107.015 ;
        RECT 63.945 104.465 69.290 105.010 ;
        RECT 69.465 104.465 74.810 105.010 ;
        RECT 74.985 104.465 80.330 105.010 ;
        RECT 80.505 104.465 85.850 105.010 ;
        RECT 86.025 104.465 88.615 105.235 ;
        RECT 89.245 104.465 89.535 105.190 ;
        RECT 91.290 105.010 91.630 105.840 ;
        RECT 93.110 105.330 93.460 106.580 ;
        RECT 96.810 105.010 97.150 105.840 ;
        RECT 98.630 105.330 98.980 106.580 ;
        RECT 102.330 105.010 102.670 105.840 ;
        RECT 104.150 105.330 104.500 106.580 ;
        RECT 107.850 105.010 108.190 105.840 ;
        RECT 109.670 105.330 110.020 106.580 ;
        RECT 111.785 105.925 114.375 107.015 ;
        RECT 111.785 105.235 112.995 105.755 ;
        RECT 113.165 105.405 114.375 105.925 ;
        RECT 115.005 105.850 115.295 107.015 ;
        RECT 115.465 106.580 120.810 107.015 ;
        RECT 120.985 106.580 126.330 107.015 ;
        RECT 126.505 106.580 131.850 107.015 ;
        RECT 132.025 106.580 137.370 107.015 ;
        RECT 89.705 104.465 95.050 105.010 ;
        RECT 95.225 104.465 100.570 105.010 ;
        RECT 100.745 104.465 106.090 105.010 ;
        RECT 106.265 104.465 111.610 105.010 ;
        RECT 111.785 104.465 114.375 105.235 ;
        RECT 115.005 104.465 115.295 105.190 ;
        RECT 117.050 105.010 117.390 105.840 ;
        RECT 118.870 105.330 119.220 106.580 ;
        RECT 122.570 105.010 122.910 105.840 ;
        RECT 124.390 105.330 124.740 106.580 ;
        RECT 128.090 105.010 128.430 105.840 ;
        RECT 129.910 105.330 130.260 106.580 ;
        RECT 133.610 105.010 133.950 105.840 ;
        RECT 135.430 105.330 135.780 106.580 ;
        RECT 138.005 105.925 139.215 107.015 ;
        RECT 138.005 105.385 138.525 105.925 ;
        RECT 138.695 105.215 139.215 105.755 ;
        RECT 115.465 104.465 120.810 105.010 ;
        RECT 120.985 104.465 126.330 105.010 ;
        RECT 126.505 104.465 131.850 105.010 ;
        RECT 132.025 104.465 137.370 105.010 ;
        RECT 138.005 104.465 139.215 105.215 ;
        RECT 50.520 104.295 139.300 104.465 ;
        RECT 50.605 103.545 51.815 104.295 ;
        RECT 52.075 103.745 52.245 104.125 ;
        RECT 52.425 103.915 52.755 104.295 ;
        RECT 52.075 103.575 52.740 103.745 ;
        RECT 52.935 103.620 53.195 104.125 ;
        RECT 53.365 103.750 58.710 104.295 ;
        RECT 50.605 103.005 51.125 103.545 ;
        RECT 51.295 102.835 51.815 103.375 ;
        RECT 52.005 103.025 52.345 103.395 ;
        RECT 52.570 103.320 52.740 103.575 ;
        RECT 52.570 102.990 52.845 103.320 ;
        RECT 52.570 102.845 52.740 102.990 ;
        RECT 50.605 101.745 51.815 102.835 ;
        RECT 52.065 102.675 52.740 102.845 ;
        RECT 53.015 102.820 53.195 103.620 ;
        RECT 54.950 102.920 55.290 103.750 ;
        RECT 59.805 103.665 60.145 104.125 ;
        RECT 60.315 103.835 60.485 104.295 ;
        RECT 60.655 103.915 61.825 104.125 ;
        RECT 60.655 103.665 60.905 103.915 ;
        RECT 61.495 103.895 61.825 103.915 ;
        RECT 62.105 103.765 62.365 104.100 ;
        RECT 62.535 103.785 62.870 104.295 ;
        RECT 63.040 103.785 63.750 104.125 ;
        RECT 59.805 103.495 60.905 103.665 ;
        RECT 61.075 103.475 61.935 103.725 ;
        RECT 52.065 101.915 52.245 102.675 ;
        RECT 52.425 101.745 52.755 102.505 ;
        RECT 52.925 101.915 53.195 102.820 ;
        RECT 56.770 102.180 57.120 103.430 ;
        RECT 59.805 103.055 60.565 103.305 ;
        RECT 60.735 103.055 61.485 103.305 ;
        RECT 61.655 102.885 61.935 103.475 ;
        RECT 53.365 101.745 58.710 102.180 ;
        RECT 59.805 101.745 60.065 102.885 ;
        RECT 60.235 102.715 61.935 102.885 ;
        RECT 60.235 101.915 60.565 102.715 ;
        RECT 60.735 101.745 60.905 102.545 ;
        RECT 61.075 101.915 61.405 102.715 ;
        RECT 61.575 101.745 61.830 102.545 ;
        RECT 62.105 102.535 62.340 103.765 ;
        RECT 62.510 102.705 62.800 103.615 ;
        RECT 62.970 103.105 63.300 103.615 ;
        RECT 63.470 103.355 63.750 103.785 ;
        RECT 63.920 103.725 64.190 104.125 ;
        RECT 64.360 103.895 64.690 104.295 ;
        RECT 64.860 103.915 66.070 104.105 ;
        RECT 64.860 103.725 65.145 103.915 ;
        RECT 66.245 103.750 71.590 104.295 ;
        RECT 63.920 103.525 65.145 103.725 ;
        RECT 65.315 103.525 66.075 103.745 ;
        RECT 63.470 103.105 64.985 103.355 ;
        RECT 65.265 103.105 65.675 103.355 ;
        RECT 63.470 102.935 63.755 103.105 ;
        RECT 65.845 102.935 66.075 103.525 ;
        RECT 63.140 102.615 63.755 102.935 ;
        RECT 63.925 102.755 66.075 102.935 ;
        RECT 67.830 102.920 68.170 103.750 ;
        RECT 71.765 103.525 75.275 104.295 ;
        RECT 76.365 103.570 76.655 104.295 ;
        RECT 76.825 103.750 82.170 104.295 ;
        RECT 82.345 103.750 87.690 104.295 ;
        RECT 87.865 103.750 93.210 104.295 ;
        RECT 93.385 103.750 98.730 104.295 ;
        RECT 63.925 102.615 65.645 102.755 ;
        RECT 62.105 101.915 62.365 102.535 ;
        RECT 62.535 101.745 62.970 102.535 ;
        RECT 63.140 101.915 63.430 102.615 ;
        RECT 63.620 102.275 65.145 102.445 ;
        RECT 63.620 101.915 63.830 102.275 ;
        RECT 64.000 101.745 64.330 102.105 ;
        RECT 64.500 102.085 65.145 102.275 ;
        RECT 65.315 102.255 65.645 102.615 ;
        RECT 65.815 102.085 66.075 102.585 ;
        RECT 69.650 102.180 70.000 103.430 ;
        RECT 71.765 103.005 73.415 103.525 ;
        RECT 73.585 102.835 75.275 103.355 ;
        RECT 78.410 102.920 78.750 103.750 ;
        RECT 64.500 101.915 66.075 102.085 ;
        RECT 66.245 101.745 71.590 102.180 ;
        RECT 71.765 101.745 75.275 102.835 ;
        RECT 76.365 101.745 76.655 102.910 ;
        RECT 80.230 102.180 80.580 103.430 ;
        RECT 83.930 102.920 84.270 103.750 ;
        RECT 85.750 102.180 86.100 103.430 ;
        RECT 89.450 102.920 89.790 103.750 ;
        RECT 91.270 102.180 91.620 103.430 ;
        RECT 94.970 102.920 95.310 103.750 ;
        RECT 98.905 103.525 101.495 104.295 ;
        RECT 102.125 103.570 102.415 104.295 ;
        RECT 102.585 103.750 107.930 104.295 ;
        RECT 108.105 103.750 113.450 104.295 ;
        RECT 113.625 103.750 118.970 104.295 ;
        RECT 119.145 103.750 124.490 104.295 ;
        RECT 96.790 102.180 97.140 103.430 ;
        RECT 98.905 103.005 100.115 103.525 ;
        RECT 100.285 102.835 101.495 103.355 ;
        RECT 104.170 102.920 104.510 103.750 ;
        RECT 76.825 101.745 82.170 102.180 ;
        RECT 82.345 101.745 87.690 102.180 ;
        RECT 87.865 101.745 93.210 102.180 ;
        RECT 93.385 101.745 98.730 102.180 ;
        RECT 98.905 101.745 101.495 102.835 ;
        RECT 102.125 101.745 102.415 102.910 ;
        RECT 105.990 102.180 106.340 103.430 ;
        RECT 109.690 102.920 110.030 103.750 ;
        RECT 111.510 102.180 111.860 103.430 ;
        RECT 115.210 102.920 115.550 103.750 ;
        RECT 117.030 102.180 117.380 103.430 ;
        RECT 120.730 102.920 121.070 103.750 ;
        RECT 124.665 103.525 127.255 104.295 ;
        RECT 127.885 103.570 128.175 104.295 ;
        RECT 128.345 103.750 133.690 104.295 ;
        RECT 122.550 102.180 122.900 103.430 ;
        RECT 124.665 103.005 125.875 103.525 ;
        RECT 126.045 102.835 127.255 103.355 ;
        RECT 129.930 102.920 130.270 103.750 ;
        RECT 133.865 103.525 137.375 104.295 ;
        RECT 138.005 103.545 139.215 104.295 ;
        RECT 102.585 101.745 107.930 102.180 ;
        RECT 108.105 101.745 113.450 102.180 ;
        RECT 113.625 101.745 118.970 102.180 ;
        RECT 119.145 101.745 124.490 102.180 ;
        RECT 124.665 101.745 127.255 102.835 ;
        RECT 127.885 101.745 128.175 102.910 ;
        RECT 131.750 102.180 132.100 103.430 ;
        RECT 133.865 103.005 135.515 103.525 ;
        RECT 135.685 102.835 137.375 103.355 ;
        RECT 128.345 101.745 133.690 102.180 ;
        RECT 133.865 101.745 137.375 102.835 ;
        RECT 138.005 102.835 138.525 103.375 ;
        RECT 138.695 103.005 139.215 103.545 ;
        RECT 138.005 101.745 139.215 102.835 ;
        RECT 50.520 101.575 139.300 101.745 ;
        RECT 50.605 100.485 51.815 101.575 ;
        RECT 50.605 99.775 51.125 100.315 ;
        RECT 51.295 99.945 51.815 100.485 ;
        RECT 52.065 100.645 52.245 101.405 ;
        RECT 52.425 100.815 52.755 101.575 ;
        RECT 52.065 100.475 52.740 100.645 ;
        RECT 52.925 100.500 53.195 101.405 ;
        RECT 53.365 101.140 58.710 101.575 ;
        RECT 52.570 100.330 52.740 100.475 ;
        RECT 52.005 99.925 52.345 100.295 ;
        RECT 52.570 100.000 52.845 100.330 ;
        RECT 50.605 99.025 51.815 99.775 ;
        RECT 52.570 99.745 52.740 100.000 ;
        RECT 52.075 99.575 52.740 99.745 ;
        RECT 53.015 99.700 53.195 100.500 ;
        RECT 52.075 99.195 52.245 99.575 ;
        RECT 52.425 99.025 52.755 99.405 ;
        RECT 52.935 99.195 53.195 99.700 ;
        RECT 54.950 99.570 55.290 100.400 ;
        RECT 56.770 99.890 57.120 101.140 ;
        RECT 58.885 100.485 62.395 101.575 ;
        RECT 58.885 99.795 60.535 100.315 ;
        RECT 60.705 99.965 62.395 100.485 ;
        RECT 63.485 100.410 63.775 101.575 ;
        RECT 63.945 101.140 69.290 101.575 ;
        RECT 69.465 101.140 74.810 101.575 ;
        RECT 74.985 101.140 80.330 101.575 ;
        RECT 80.505 101.140 85.850 101.575 ;
        RECT 53.365 99.025 58.710 99.570 ;
        RECT 58.885 99.025 62.395 99.795 ;
        RECT 63.485 99.025 63.775 99.750 ;
        RECT 65.530 99.570 65.870 100.400 ;
        RECT 67.350 99.890 67.700 101.140 ;
        RECT 71.050 99.570 71.390 100.400 ;
        RECT 72.870 99.890 73.220 101.140 ;
        RECT 76.570 99.570 76.910 100.400 ;
        RECT 78.390 99.890 78.740 101.140 ;
        RECT 82.090 99.570 82.430 100.400 ;
        RECT 83.910 99.890 84.260 101.140 ;
        RECT 86.025 100.485 88.615 101.575 ;
        RECT 86.025 99.795 87.235 100.315 ;
        RECT 87.405 99.965 88.615 100.485 ;
        RECT 89.245 100.410 89.535 101.575 ;
        RECT 89.705 101.140 95.050 101.575 ;
        RECT 95.225 101.140 100.570 101.575 ;
        RECT 100.745 101.140 106.090 101.575 ;
        RECT 106.265 101.140 111.610 101.575 ;
        RECT 63.945 99.025 69.290 99.570 ;
        RECT 69.465 99.025 74.810 99.570 ;
        RECT 74.985 99.025 80.330 99.570 ;
        RECT 80.505 99.025 85.850 99.570 ;
        RECT 86.025 99.025 88.615 99.795 ;
        RECT 89.245 99.025 89.535 99.750 ;
        RECT 91.290 99.570 91.630 100.400 ;
        RECT 93.110 99.890 93.460 101.140 ;
        RECT 96.810 99.570 97.150 100.400 ;
        RECT 98.630 99.890 98.980 101.140 ;
        RECT 102.330 99.570 102.670 100.400 ;
        RECT 104.150 99.890 104.500 101.140 ;
        RECT 107.850 99.570 108.190 100.400 ;
        RECT 109.670 99.890 110.020 101.140 ;
        RECT 111.785 100.485 114.375 101.575 ;
        RECT 111.785 99.795 112.995 100.315 ;
        RECT 113.165 99.965 114.375 100.485 ;
        RECT 115.005 100.410 115.295 101.575 ;
        RECT 115.465 101.140 120.810 101.575 ;
        RECT 120.985 101.140 126.330 101.575 ;
        RECT 126.505 101.140 131.850 101.575 ;
        RECT 132.025 101.140 137.370 101.575 ;
        RECT 89.705 99.025 95.050 99.570 ;
        RECT 95.225 99.025 100.570 99.570 ;
        RECT 100.745 99.025 106.090 99.570 ;
        RECT 106.265 99.025 111.610 99.570 ;
        RECT 111.785 99.025 114.375 99.795 ;
        RECT 115.005 99.025 115.295 99.750 ;
        RECT 117.050 99.570 117.390 100.400 ;
        RECT 118.870 99.890 119.220 101.140 ;
        RECT 122.570 99.570 122.910 100.400 ;
        RECT 124.390 99.890 124.740 101.140 ;
        RECT 128.090 99.570 128.430 100.400 ;
        RECT 129.910 99.890 130.260 101.140 ;
        RECT 133.610 99.570 133.950 100.400 ;
        RECT 135.430 99.890 135.780 101.140 ;
        RECT 138.005 100.485 139.215 101.575 ;
        RECT 138.005 99.945 138.525 100.485 ;
        RECT 138.695 99.775 139.215 100.315 ;
        RECT 115.465 99.025 120.810 99.570 ;
        RECT 120.985 99.025 126.330 99.570 ;
        RECT 126.505 99.025 131.850 99.570 ;
        RECT 132.025 99.025 137.370 99.570 ;
        RECT 138.005 99.025 139.215 99.775 ;
        RECT 50.520 98.855 139.300 99.025 ;
        RECT 50.605 98.105 51.815 98.855 ;
        RECT 51.985 98.310 57.330 98.855 ;
        RECT 50.605 97.565 51.125 98.105 ;
        RECT 51.295 97.395 51.815 97.935 ;
        RECT 53.570 97.480 53.910 98.310 ;
        RECT 57.505 98.085 60.095 98.855 ;
        RECT 60.815 98.305 60.985 98.685 ;
        RECT 61.165 98.475 61.495 98.855 ;
        RECT 60.815 98.135 61.480 98.305 ;
        RECT 61.675 98.180 61.935 98.685 ;
        RECT 62.105 98.310 67.450 98.855 ;
        RECT 67.625 98.310 72.970 98.855 ;
        RECT 50.605 96.305 51.815 97.395 ;
        RECT 55.390 96.740 55.740 97.990 ;
        RECT 57.505 97.565 58.715 98.085 ;
        RECT 58.885 97.395 60.095 97.915 ;
        RECT 60.745 97.585 61.075 97.955 ;
        RECT 61.310 97.880 61.480 98.135 ;
        RECT 61.310 97.550 61.595 97.880 ;
        RECT 61.310 97.405 61.480 97.550 ;
        RECT 51.985 96.305 57.330 96.740 ;
        RECT 57.505 96.305 60.095 97.395 ;
        RECT 60.815 97.235 61.480 97.405 ;
        RECT 61.765 97.380 61.935 98.180 ;
        RECT 63.690 97.480 64.030 98.310 ;
        RECT 60.815 96.475 60.985 97.235 ;
        RECT 61.165 96.305 61.495 97.065 ;
        RECT 61.665 96.475 61.935 97.380 ;
        RECT 65.510 96.740 65.860 97.990 ;
        RECT 69.210 97.480 69.550 98.310 ;
        RECT 73.145 98.085 75.735 98.855 ;
        RECT 76.365 98.130 76.655 98.855 ;
        RECT 76.825 98.310 82.170 98.855 ;
        RECT 82.345 98.310 87.690 98.855 ;
        RECT 87.865 98.310 93.210 98.855 ;
        RECT 93.385 98.310 98.730 98.855 ;
        RECT 71.030 96.740 71.380 97.990 ;
        RECT 73.145 97.565 74.355 98.085 ;
        RECT 74.525 97.395 75.735 97.915 ;
        RECT 78.410 97.480 78.750 98.310 ;
        RECT 62.105 96.305 67.450 96.740 ;
        RECT 67.625 96.305 72.970 96.740 ;
        RECT 73.145 96.305 75.735 97.395 ;
        RECT 76.365 96.305 76.655 97.470 ;
        RECT 80.230 96.740 80.580 97.990 ;
        RECT 83.930 97.480 84.270 98.310 ;
        RECT 85.750 96.740 86.100 97.990 ;
        RECT 89.450 97.480 89.790 98.310 ;
        RECT 91.270 96.740 91.620 97.990 ;
        RECT 94.970 97.480 95.310 98.310 ;
        RECT 98.905 98.085 101.495 98.855 ;
        RECT 102.125 98.130 102.415 98.855 ;
        RECT 102.585 98.310 107.930 98.855 ;
        RECT 108.105 98.310 113.450 98.855 ;
        RECT 113.625 98.310 118.970 98.855 ;
        RECT 119.145 98.310 124.490 98.855 ;
        RECT 96.790 96.740 97.140 97.990 ;
        RECT 98.905 97.565 100.115 98.085 ;
        RECT 100.285 97.395 101.495 97.915 ;
        RECT 104.170 97.480 104.510 98.310 ;
        RECT 76.825 96.305 82.170 96.740 ;
        RECT 82.345 96.305 87.690 96.740 ;
        RECT 87.865 96.305 93.210 96.740 ;
        RECT 93.385 96.305 98.730 96.740 ;
        RECT 98.905 96.305 101.495 97.395 ;
        RECT 102.125 96.305 102.415 97.470 ;
        RECT 105.990 96.740 106.340 97.990 ;
        RECT 109.690 97.480 110.030 98.310 ;
        RECT 111.510 96.740 111.860 97.990 ;
        RECT 115.210 97.480 115.550 98.310 ;
        RECT 117.030 96.740 117.380 97.990 ;
        RECT 120.730 97.480 121.070 98.310 ;
        RECT 124.665 98.085 127.255 98.855 ;
        RECT 127.885 98.130 128.175 98.855 ;
        RECT 128.345 98.310 133.690 98.855 ;
        RECT 122.550 96.740 122.900 97.990 ;
        RECT 124.665 97.565 125.875 98.085 ;
        RECT 126.045 97.395 127.255 97.915 ;
        RECT 129.930 97.480 130.270 98.310 ;
        RECT 133.865 98.085 137.375 98.855 ;
        RECT 138.005 98.105 139.215 98.855 ;
        RECT 102.585 96.305 107.930 96.740 ;
        RECT 108.105 96.305 113.450 96.740 ;
        RECT 113.625 96.305 118.970 96.740 ;
        RECT 119.145 96.305 124.490 96.740 ;
        RECT 124.665 96.305 127.255 97.395 ;
        RECT 127.885 96.305 128.175 97.470 ;
        RECT 131.750 96.740 132.100 97.990 ;
        RECT 133.865 97.565 135.515 98.085 ;
        RECT 135.685 97.395 137.375 97.915 ;
        RECT 128.345 96.305 133.690 96.740 ;
        RECT 133.865 96.305 137.375 97.395 ;
        RECT 138.005 97.395 138.525 97.935 ;
        RECT 138.695 97.565 139.215 98.105 ;
        RECT 138.005 96.305 139.215 97.395 ;
        RECT 50.520 96.135 139.300 96.305 ;
        RECT 50.605 95.045 51.815 96.135 ;
        RECT 51.985 95.700 57.330 96.135 ;
        RECT 50.605 94.335 51.125 94.875 ;
        RECT 51.295 94.505 51.815 95.045 ;
        RECT 50.605 93.585 51.815 94.335 ;
        RECT 53.570 94.130 53.910 94.960 ;
        RECT 55.390 94.450 55.740 95.700 ;
        RECT 57.505 95.045 61.015 96.135 ;
        RECT 57.505 94.355 59.155 94.875 ;
        RECT 59.325 94.525 61.015 95.045 ;
        RECT 61.645 94.995 61.905 96.135 ;
        RECT 62.075 94.985 62.405 95.965 ;
        RECT 62.575 94.995 62.855 96.135 ;
        RECT 61.665 94.575 62.000 94.825 ;
        RECT 62.170 94.385 62.340 94.985 ;
        RECT 63.485 94.970 63.775 96.135 ;
        RECT 63.945 95.700 69.290 96.135 ;
        RECT 69.465 95.700 74.810 96.135 ;
        RECT 74.985 95.700 80.330 96.135 ;
        RECT 80.505 95.700 85.850 96.135 ;
        RECT 62.510 94.555 62.845 94.825 ;
        RECT 51.985 93.585 57.330 94.130 ;
        RECT 57.505 93.585 61.015 94.355 ;
        RECT 61.645 93.755 62.340 94.385 ;
        RECT 62.545 93.585 62.855 94.385 ;
        RECT 63.485 93.585 63.775 94.310 ;
        RECT 65.530 94.130 65.870 94.960 ;
        RECT 67.350 94.450 67.700 95.700 ;
        RECT 71.050 94.130 71.390 94.960 ;
        RECT 72.870 94.450 73.220 95.700 ;
        RECT 76.570 94.130 76.910 94.960 ;
        RECT 78.390 94.450 78.740 95.700 ;
        RECT 82.090 94.130 82.430 94.960 ;
        RECT 83.910 94.450 84.260 95.700 ;
        RECT 86.025 95.045 88.615 96.135 ;
        RECT 86.025 94.355 87.235 94.875 ;
        RECT 87.405 94.525 88.615 95.045 ;
        RECT 89.245 94.970 89.535 96.135 ;
        RECT 89.705 95.700 95.050 96.135 ;
        RECT 95.225 95.700 100.570 96.135 ;
        RECT 100.745 95.700 106.090 96.135 ;
        RECT 106.265 95.700 111.610 96.135 ;
        RECT 63.945 93.585 69.290 94.130 ;
        RECT 69.465 93.585 74.810 94.130 ;
        RECT 74.985 93.585 80.330 94.130 ;
        RECT 80.505 93.585 85.850 94.130 ;
        RECT 86.025 93.585 88.615 94.355 ;
        RECT 89.245 93.585 89.535 94.310 ;
        RECT 91.290 94.130 91.630 94.960 ;
        RECT 93.110 94.450 93.460 95.700 ;
        RECT 96.810 94.130 97.150 94.960 ;
        RECT 98.630 94.450 98.980 95.700 ;
        RECT 102.330 94.130 102.670 94.960 ;
        RECT 104.150 94.450 104.500 95.700 ;
        RECT 107.850 94.130 108.190 94.960 ;
        RECT 109.670 94.450 110.020 95.700 ;
        RECT 111.785 95.045 114.375 96.135 ;
        RECT 111.785 94.355 112.995 94.875 ;
        RECT 113.165 94.525 114.375 95.045 ;
        RECT 115.005 94.970 115.295 96.135 ;
        RECT 115.465 95.700 120.810 96.135 ;
        RECT 120.985 95.700 126.330 96.135 ;
        RECT 126.505 95.700 131.850 96.135 ;
        RECT 132.025 95.700 137.370 96.135 ;
        RECT 89.705 93.585 95.050 94.130 ;
        RECT 95.225 93.585 100.570 94.130 ;
        RECT 100.745 93.585 106.090 94.130 ;
        RECT 106.265 93.585 111.610 94.130 ;
        RECT 111.785 93.585 114.375 94.355 ;
        RECT 115.005 93.585 115.295 94.310 ;
        RECT 117.050 94.130 117.390 94.960 ;
        RECT 118.870 94.450 119.220 95.700 ;
        RECT 122.570 94.130 122.910 94.960 ;
        RECT 124.390 94.450 124.740 95.700 ;
        RECT 128.090 94.130 128.430 94.960 ;
        RECT 129.910 94.450 130.260 95.700 ;
        RECT 133.610 94.130 133.950 94.960 ;
        RECT 135.430 94.450 135.780 95.700 ;
        RECT 138.005 95.045 139.215 96.135 ;
        RECT 138.005 94.505 138.525 95.045 ;
        RECT 138.695 94.335 139.215 94.875 ;
        RECT 115.465 93.585 120.810 94.130 ;
        RECT 120.985 93.585 126.330 94.130 ;
        RECT 126.505 93.585 131.850 94.130 ;
        RECT 132.025 93.585 137.370 94.130 ;
        RECT 138.005 93.585 139.215 94.335 ;
        RECT 50.520 93.415 139.300 93.585 ;
        RECT 50.605 92.665 51.815 93.415 ;
        RECT 50.605 92.125 51.125 92.665 ;
        RECT 51.985 92.645 55.495 93.415 ;
        RECT 51.295 91.955 51.815 92.495 ;
        RECT 51.985 92.125 53.635 92.645 ;
        RECT 56.860 92.605 57.105 93.210 ;
        RECT 57.325 92.880 57.835 93.415 ;
        RECT 53.805 91.955 55.495 92.475 ;
        RECT 50.605 90.865 51.815 91.955 ;
        RECT 51.985 90.865 55.495 91.955 ;
        RECT 56.585 92.435 57.815 92.605 ;
        RECT 56.585 91.625 56.925 92.435 ;
        RECT 57.095 91.870 57.845 92.060 ;
        RECT 56.585 91.215 57.100 91.625 ;
        RECT 57.335 90.865 57.505 91.625 ;
        RECT 57.675 91.205 57.845 91.870 ;
        RECT 58.015 91.885 58.205 93.245 ;
        RECT 58.375 93.075 58.650 93.245 ;
        RECT 58.375 92.905 58.655 93.075 ;
        RECT 58.375 92.085 58.650 92.905 ;
        RECT 58.840 92.880 59.370 93.245 ;
        RECT 59.795 93.015 60.125 93.415 ;
        RECT 59.195 92.845 59.370 92.880 ;
        RECT 58.855 91.885 59.025 92.685 ;
        RECT 58.015 91.715 59.025 91.885 ;
        RECT 59.195 92.675 60.125 92.845 ;
        RECT 60.295 92.675 60.550 93.245 ;
        RECT 59.195 91.545 59.365 92.675 ;
        RECT 59.955 92.505 60.125 92.675 ;
        RECT 58.240 91.375 59.365 91.545 ;
        RECT 59.535 92.175 59.730 92.505 ;
        RECT 59.955 92.175 60.210 92.505 ;
        RECT 59.535 91.205 59.705 92.175 ;
        RECT 60.380 92.005 60.550 92.675 ;
        RECT 57.675 91.035 59.705 91.205 ;
        RECT 59.875 90.865 60.045 92.005 ;
        RECT 60.215 91.035 60.550 92.005 ;
        RECT 60.730 92.675 60.985 93.245 ;
        RECT 61.155 93.015 61.485 93.415 ;
        RECT 61.910 92.880 62.440 93.245 ;
        RECT 61.910 92.845 62.085 92.880 ;
        RECT 61.155 92.675 62.085 92.845 ;
        RECT 60.730 92.005 60.900 92.675 ;
        RECT 61.155 92.505 61.325 92.675 ;
        RECT 61.070 92.175 61.325 92.505 ;
        RECT 61.550 92.175 61.745 92.505 ;
        RECT 60.730 91.035 61.065 92.005 ;
        RECT 61.235 90.865 61.405 92.005 ;
        RECT 61.575 91.205 61.745 92.175 ;
        RECT 61.915 91.545 62.085 92.675 ;
        RECT 62.255 91.885 62.425 92.685 ;
        RECT 62.630 92.395 62.905 93.245 ;
        RECT 62.625 92.225 62.905 92.395 ;
        RECT 62.630 92.085 62.905 92.225 ;
        RECT 63.075 91.885 63.265 93.245 ;
        RECT 63.445 92.880 63.955 93.415 ;
        RECT 64.175 92.605 64.420 93.210 ;
        RECT 63.465 92.435 64.695 92.605 ;
        RECT 64.905 92.595 65.135 93.415 ;
        RECT 65.305 92.615 65.635 93.245 ;
        RECT 62.255 91.715 63.265 91.885 ;
        RECT 63.435 91.870 64.185 92.060 ;
        RECT 61.915 91.375 63.040 91.545 ;
        RECT 63.435 91.205 63.605 91.870 ;
        RECT 64.355 91.625 64.695 92.435 ;
        RECT 64.885 92.175 65.215 92.425 ;
        RECT 65.385 92.015 65.635 92.615 ;
        RECT 65.805 92.595 66.015 93.415 ;
        RECT 66.285 92.595 66.515 93.415 ;
        RECT 66.685 92.615 67.015 93.245 ;
        RECT 66.265 92.175 66.595 92.425 ;
        RECT 66.765 92.015 67.015 92.615 ;
        RECT 67.185 92.595 67.395 93.415 ;
        RECT 67.625 92.870 72.970 93.415 ;
        RECT 69.210 92.040 69.550 92.870 ;
        RECT 73.145 92.645 75.735 93.415 ;
        RECT 76.365 92.690 76.655 93.415 ;
        RECT 76.825 92.870 82.170 93.415 ;
        RECT 82.345 92.870 87.690 93.415 ;
        RECT 87.865 92.870 93.210 93.415 ;
        RECT 93.385 92.870 98.730 93.415 ;
        RECT 61.575 91.035 63.605 91.205 ;
        RECT 63.775 90.865 63.945 91.625 ;
        RECT 64.180 91.215 64.695 91.625 ;
        RECT 64.905 90.865 65.135 92.005 ;
        RECT 65.305 91.035 65.635 92.015 ;
        RECT 65.805 90.865 66.015 92.005 ;
        RECT 66.285 90.865 66.515 92.005 ;
        RECT 66.685 91.035 67.015 92.015 ;
        RECT 67.185 90.865 67.395 92.005 ;
        RECT 71.030 91.300 71.380 92.550 ;
        RECT 73.145 92.125 74.355 92.645 ;
        RECT 74.525 91.955 75.735 92.475 ;
        RECT 78.410 92.040 78.750 92.870 ;
        RECT 67.625 90.865 72.970 91.300 ;
        RECT 73.145 90.865 75.735 91.955 ;
        RECT 76.365 90.865 76.655 92.030 ;
        RECT 80.230 91.300 80.580 92.550 ;
        RECT 83.930 92.040 84.270 92.870 ;
        RECT 85.750 91.300 86.100 92.550 ;
        RECT 89.450 92.040 89.790 92.870 ;
        RECT 91.270 91.300 91.620 92.550 ;
        RECT 94.970 92.040 95.310 92.870 ;
        RECT 98.905 92.645 101.495 93.415 ;
        RECT 102.125 92.690 102.415 93.415 ;
        RECT 102.585 92.870 107.930 93.415 ;
        RECT 108.105 92.870 113.450 93.415 ;
        RECT 113.625 92.870 118.970 93.415 ;
        RECT 119.145 92.870 124.490 93.415 ;
        RECT 96.790 91.300 97.140 92.550 ;
        RECT 98.905 92.125 100.115 92.645 ;
        RECT 100.285 91.955 101.495 92.475 ;
        RECT 104.170 92.040 104.510 92.870 ;
        RECT 76.825 90.865 82.170 91.300 ;
        RECT 82.345 90.865 87.690 91.300 ;
        RECT 87.865 90.865 93.210 91.300 ;
        RECT 93.385 90.865 98.730 91.300 ;
        RECT 98.905 90.865 101.495 91.955 ;
        RECT 102.125 90.865 102.415 92.030 ;
        RECT 105.990 91.300 106.340 92.550 ;
        RECT 109.690 92.040 110.030 92.870 ;
        RECT 111.510 91.300 111.860 92.550 ;
        RECT 115.210 92.040 115.550 92.870 ;
        RECT 117.030 91.300 117.380 92.550 ;
        RECT 120.730 92.040 121.070 92.870 ;
        RECT 124.665 92.645 127.255 93.415 ;
        RECT 127.885 92.690 128.175 93.415 ;
        RECT 128.345 92.870 133.690 93.415 ;
        RECT 122.550 91.300 122.900 92.550 ;
        RECT 124.665 92.125 125.875 92.645 ;
        RECT 126.045 91.955 127.255 92.475 ;
        RECT 129.930 92.040 130.270 92.870 ;
        RECT 133.865 92.645 137.375 93.415 ;
        RECT 138.005 92.665 139.215 93.415 ;
        RECT 102.585 90.865 107.930 91.300 ;
        RECT 108.105 90.865 113.450 91.300 ;
        RECT 113.625 90.865 118.970 91.300 ;
        RECT 119.145 90.865 124.490 91.300 ;
        RECT 124.665 90.865 127.255 91.955 ;
        RECT 127.885 90.865 128.175 92.030 ;
        RECT 131.750 91.300 132.100 92.550 ;
        RECT 133.865 92.125 135.515 92.645 ;
        RECT 135.685 91.955 137.375 92.475 ;
        RECT 128.345 90.865 133.690 91.300 ;
        RECT 133.865 90.865 137.375 91.955 ;
        RECT 138.005 91.955 138.525 92.495 ;
        RECT 138.695 92.125 139.215 92.665 ;
        RECT 138.005 90.865 139.215 91.955 ;
        RECT 50.520 90.695 139.300 90.865 ;
        RECT 50.605 89.605 51.815 90.695 ;
        RECT 51.985 90.260 57.330 90.695 ;
        RECT 50.605 88.895 51.125 89.435 ;
        RECT 51.295 89.065 51.815 89.605 ;
        RECT 50.605 88.145 51.815 88.895 ;
        RECT 53.570 88.690 53.910 89.520 ;
        RECT 55.390 89.010 55.740 90.260 ;
        RECT 57.505 89.605 60.095 90.695 ;
        RECT 57.505 88.915 58.715 89.435 ;
        RECT 58.885 89.085 60.095 89.605 ;
        RECT 60.345 89.765 60.525 90.525 ;
        RECT 60.705 89.935 61.035 90.695 ;
        RECT 60.345 89.595 61.020 89.765 ;
        RECT 61.205 89.620 61.475 90.525 ;
        RECT 60.850 89.450 61.020 89.595 ;
        RECT 60.285 89.045 60.625 89.415 ;
        RECT 60.850 89.120 61.125 89.450 ;
        RECT 51.985 88.145 57.330 88.690 ;
        RECT 57.505 88.145 60.095 88.915 ;
        RECT 60.850 88.865 61.020 89.120 ;
        RECT 60.355 88.695 61.020 88.865 ;
        RECT 61.295 88.820 61.475 89.620 ;
        RECT 61.685 89.555 61.915 90.695 ;
        RECT 62.085 89.545 62.415 90.525 ;
        RECT 62.585 89.555 62.795 90.695 ;
        RECT 61.665 89.135 61.995 89.385 ;
        RECT 60.355 88.315 60.525 88.695 ;
        RECT 60.705 88.145 61.035 88.525 ;
        RECT 61.215 88.315 61.475 88.820 ;
        RECT 61.685 88.145 61.915 88.965 ;
        RECT 62.165 88.945 62.415 89.545 ;
        RECT 63.485 89.530 63.775 90.695 ;
        RECT 63.945 90.260 69.290 90.695 ;
        RECT 69.465 90.260 74.810 90.695 ;
        RECT 74.985 90.260 80.330 90.695 ;
        RECT 80.505 90.260 85.850 90.695 ;
        RECT 62.085 88.315 62.415 88.945 ;
        RECT 62.585 88.145 62.795 88.965 ;
        RECT 63.485 88.145 63.775 88.870 ;
        RECT 65.530 88.690 65.870 89.520 ;
        RECT 67.350 89.010 67.700 90.260 ;
        RECT 71.050 88.690 71.390 89.520 ;
        RECT 72.870 89.010 73.220 90.260 ;
        RECT 76.570 88.690 76.910 89.520 ;
        RECT 78.390 89.010 78.740 90.260 ;
        RECT 82.090 88.690 82.430 89.520 ;
        RECT 83.910 89.010 84.260 90.260 ;
        RECT 86.025 89.605 88.615 90.695 ;
        RECT 86.025 88.915 87.235 89.435 ;
        RECT 87.405 89.085 88.615 89.605 ;
        RECT 89.245 89.530 89.535 90.695 ;
        RECT 89.705 90.260 95.050 90.695 ;
        RECT 95.225 90.260 100.570 90.695 ;
        RECT 100.745 90.260 106.090 90.695 ;
        RECT 106.265 90.260 111.610 90.695 ;
        RECT 63.945 88.145 69.290 88.690 ;
        RECT 69.465 88.145 74.810 88.690 ;
        RECT 74.985 88.145 80.330 88.690 ;
        RECT 80.505 88.145 85.850 88.690 ;
        RECT 86.025 88.145 88.615 88.915 ;
        RECT 89.245 88.145 89.535 88.870 ;
        RECT 91.290 88.690 91.630 89.520 ;
        RECT 93.110 89.010 93.460 90.260 ;
        RECT 96.810 88.690 97.150 89.520 ;
        RECT 98.630 89.010 98.980 90.260 ;
        RECT 102.330 88.690 102.670 89.520 ;
        RECT 104.150 89.010 104.500 90.260 ;
        RECT 107.850 88.690 108.190 89.520 ;
        RECT 109.670 89.010 110.020 90.260 ;
        RECT 111.785 89.605 114.375 90.695 ;
        RECT 111.785 88.915 112.995 89.435 ;
        RECT 113.165 89.085 114.375 89.605 ;
        RECT 115.005 89.530 115.295 90.695 ;
        RECT 115.465 90.260 120.810 90.695 ;
        RECT 120.985 90.260 126.330 90.695 ;
        RECT 126.505 90.260 131.850 90.695 ;
        RECT 132.025 90.260 137.370 90.695 ;
        RECT 89.705 88.145 95.050 88.690 ;
        RECT 95.225 88.145 100.570 88.690 ;
        RECT 100.745 88.145 106.090 88.690 ;
        RECT 106.265 88.145 111.610 88.690 ;
        RECT 111.785 88.145 114.375 88.915 ;
        RECT 115.005 88.145 115.295 88.870 ;
        RECT 117.050 88.690 117.390 89.520 ;
        RECT 118.870 89.010 119.220 90.260 ;
        RECT 122.570 88.690 122.910 89.520 ;
        RECT 124.390 89.010 124.740 90.260 ;
        RECT 128.090 88.690 128.430 89.520 ;
        RECT 129.910 89.010 130.260 90.260 ;
        RECT 133.610 88.690 133.950 89.520 ;
        RECT 135.430 89.010 135.780 90.260 ;
        RECT 138.005 89.605 139.215 90.695 ;
        RECT 138.005 89.065 138.525 89.605 ;
        RECT 138.695 88.895 139.215 89.435 ;
        RECT 115.465 88.145 120.810 88.690 ;
        RECT 120.985 88.145 126.330 88.690 ;
        RECT 126.505 88.145 131.850 88.690 ;
        RECT 132.025 88.145 137.370 88.690 ;
        RECT 138.005 88.145 139.215 88.895 ;
        RECT 50.520 87.975 139.300 88.145 ;
        RECT 50.605 87.225 51.815 87.975 ;
        RECT 51.985 87.430 57.330 87.975 ;
        RECT 57.505 87.430 62.850 87.975 ;
        RECT 63.025 87.430 68.370 87.975 ;
        RECT 68.545 87.430 73.890 87.975 ;
        RECT 50.605 86.685 51.125 87.225 ;
        RECT 51.295 86.515 51.815 87.055 ;
        RECT 53.570 86.600 53.910 87.430 ;
        RECT 50.605 85.425 51.815 86.515 ;
        RECT 55.390 85.860 55.740 87.110 ;
        RECT 59.090 86.600 59.430 87.430 ;
        RECT 60.910 85.860 61.260 87.110 ;
        RECT 64.610 86.600 64.950 87.430 ;
        RECT 66.430 85.860 66.780 87.110 ;
        RECT 70.130 86.600 70.470 87.430 ;
        RECT 74.065 87.205 75.735 87.975 ;
        RECT 76.365 87.250 76.655 87.975 ;
        RECT 76.825 87.430 82.170 87.975 ;
        RECT 82.345 87.430 87.690 87.975 ;
        RECT 87.865 87.430 93.210 87.975 ;
        RECT 93.385 87.430 98.730 87.975 ;
        RECT 71.950 85.860 72.300 87.110 ;
        RECT 74.065 86.685 74.815 87.205 ;
        RECT 74.985 86.515 75.735 87.035 ;
        RECT 78.410 86.600 78.750 87.430 ;
        RECT 51.985 85.425 57.330 85.860 ;
        RECT 57.505 85.425 62.850 85.860 ;
        RECT 63.025 85.425 68.370 85.860 ;
        RECT 68.545 85.425 73.890 85.860 ;
        RECT 74.065 85.425 75.735 86.515 ;
        RECT 76.365 85.425 76.655 86.590 ;
        RECT 80.230 85.860 80.580 87.110 ;
        RECT 83.930 86.600 84.270 87.430 ;
        RECT 85.750 85.860 86.100 87.110 ;
        RECT 89.450 86.600 89.790 87.430 ;
        RECT 91.270 85.860 91.620 87.110 ;
        RECT 94.970 86.600 95.310 87.430 ;
        RECT 98.905 87.205 101.495 87.975 ;
        RECT 102.125 87.250 102.415 87.975 ;
        RECT 102.585 87.430 107.930 87.975 ;
        RECT 108.105 87.430 113.450 87.975 ;
        RECT 113.625 87.430 118.970 87.975 ;
        RECT 119.145 87.430 124.490 87.975 ;
        RECT 96.790 85.860 97.140 87.110 ;
        RECT 98.905 86.685 100.115 87.205 ;
        RECT 100.285 86.515 101.495 87.035 ;
        RECT 104.170 86.600 104.510 87.430 ;
        RECT 76.825 85.425 82.170 85.860 ;
        RECT 82.345 85.425 87.690 85.860 ;
        RECT 87.865 85.425 93.210 85.860 ;
        RECT 93.385 85.425 98.730 85.860 ;
        RECT 98.905 85.425 101.495 86.515 ;
        RECT 102.125 85.425 102.415 86.590 ;
        RECT 105.990 85.860 106.340 87.110 ;
        RECT 109.690 86.600 110.030 87.430 ;
        RECT 111.510 85.860 111.860 87.110 ;
        RECT 115.210 86.600 115.550 87.430 ;
        RECT 117.030 85.860 117.380 87.110 ;
        RECT 120.730 86.600 121.070 87.430 ;
        RECT 124.665 87.205 127.255 87.975 ;
        RECT 127.885 87.250 128.175 87.975 ;
        RECT 128.345 87.430 133.690 87.975 ;
        RECT 122.550 85.860 122.900 87.110 ;
        RECT 124.665 86.685 125.875 87.205 ;
        RECT 126.045 86.515 127.255 87.035 ;
        RECT 129.930 86.600 130.270 87.430 ;
        RECT 133.865 87.205 137.375 87.975 ;
        RECT 138.005 87.225 139.215 87.975 ;
        RECT 102.585 85.425 107.930 85.860 ;
        RECT 108.105 85.425 113.450 85.860 ;
        RECT 113.625 85.425 118.970 85.860 ;
        RECT 119.145 85.425 124.490 85.860 ;
        RECT 124.665 85.425 127.255 86.515 ;
        RECT 127.885 85.425 128.175 86.590 ;
        RECT 131.750 85.860 132.100 87.110 ;
        RECT 133.865 86.685 135.515 87.205 ;
        RECT 135.685 86.515 137.375 87.035 ;
        RECT 128.345 85.425 133.690 85.860 ;
        RECT 133.865 85.425 137.375 86.515 ;
        RECT 138.005 86.515 138.525 87.055 ;
        RECT 138.695 86.685 139.215 87.225 ;
        RECT 138.005 85.425 139.215 86.515 ;
        RECT 50.520 85.255 139.300 85.425 ;
        RECT 50.605 84.165 51.815 85.255 ;
        RECT 51.985 84.820 57.330 85.255 ;
        RECT 57.505 84.820 62.850 85.255 ;
        RECT 50.605 83.455 51.125 83.995 ;
        RECT 51.295 83.625 51.815 84.165 ;
        RECT 50.605 82.705 51.815 83.455 ;
        RECT 53.570 83.250 53.910 84.080 ;
        RECT 55.390 83.570 55.740 84.820 ;
        RECT 59.090 83.250 59.430 84.080 ;
        RECT 60.910 83.570 61.260 84.820 ;
        RECT 63.485 84.090 63.775 85.255 ;
        RECT 63.945 84.820 69.290 85.255 ;
        RECT 69.465 84.820 74.810 85.255 ;
        RECT 74.985 84.820 80.330 85.255 ;
        RECT 80.505 84.820 85.850 85.255 ;
        RECT 51.985 82.705 57.330 83.250 ;
        RECT 57.505 82.705 62.850 83.250 ;
        RECT 63.485 82.705 63.775 83.430 ;
        RECT 65.530 83.250 65.870 84.080 ;
        RECT 67.350 83.570 67.700 84.820 ;
        RECT 71.050 83.250 71.390 84.080 ;
        RECT 72.870 83.570 73.220 84.820 ;
        RECT 76.570 83.250 76.910 84.080 ;
        RECT 78.390 83.570 78.740 84.820 ;
        RECT 82.090 83.250 82.430 84.080 ;
        RECT 83.910 83.570 84.260 84.820 ;
        RECT 86.025 84.165 88.615 85.255 ;
        RECT 86.025 83.475 87.235 83.995 ;
        RECT 87.405 83.645 88.615 84.165 ;
        RECT 89.245 84.090 89.535 85.255 ;
        RECT 89.705 84.820 95.050 85.255 ;
        RECT 95.225 84.820 100.570 85.255 ;
        RECT 100.745 84.820 106.090 85.255 ;
        RECT 106.265 84.820 111.610 85.255 ;
        RECT 63.945 82.705 69.290 83.250 ;
        RECT 69.465 82.705 74.810 83.250 ;
        RECT 74.985 82.705 80.330 83.250 ;
        RECT 80.505 82.705 85.850 83.250 ;
        RECT 86.025 82.705 88.615 83.475 ;
        RECT 89.245 82.705 89.535 83.430 ;
        RECT 91.290 83.250 91.630 84.080 ;
        RECT 93.110 83.570 93.460 84.820 ;
        RECT 96.810 83.250 97.150 84.080 ;
        RECT 98.630 83.570 98.980 84.820 ;
        RECT 102.330 83.250 102.670 84.080 ;
        RECT 104.150 83.570 104.500 84.820 ;
        RECT 107.850 83.250 108.190 84.080 ;
        RECT 109.670 83.570 110.020 84.820 ;
        RECT 111.785 84.165 114.375 85.255 ;
        RECT 111.785 83.475 112.995 83.995 ;
        RECT 113.165 83.645 114.375 84.165 ;
        RECT 115.005 84.090 115.295 85.255 ;
        RECT 115.465 84.820 120.810 85.255 ;
        RECT 120.985 84.820 126.330 85.255 ;
        RECT 126.505 84.820 131.850 85.255 ;
        RECT 132.025 84.820 137.370 85.255 ;
        RECT 89.705 82.705 95.050 83.250 ;
        RECT 95.225 82.705 100.570 83.250 ;
        RECT 100.745 82.705 106.090 83.250 ;
        RECT 106.265 82.705 111.610 83.250 ;
        RECT 111.785 82.705 114.375 83.475 ;
        RECT 115.005 82.705 115.295 83.430 ;
        RECT 117.050 83.250 117.390 84.080 ;
        RECT 118.870 83.570 119.220 84.820 ;
        RECT 122.570 83.250 122.910 84.080 ;
        RECT 124.390 83.570 124.740 84.820 ;
        RECT 128.090 83.250 128.430 84.080 ;
        RECT 129.910 83.570 130.260 84.820 ;
        RECT 133.610 83.250 133.950 84.080 ;
        RECT 135.430 83.570 135.780 84.820 ;
        RECT 138.005 84.165 139.215 85.255 ;
        RECT 138.005 83.625 138.525 84.165 ;
        RECT 138.695 83.455 139.215 83.995 ;
        RECT 115.465 82.705 120.810 83.250 ;
        RECT 120.985 82.705 126.330 83.250 ;
        RECT 126.505 82.705 131.850 83.250 ;
        RECT 132.025 82.705 137.370 83.250 ;
        RECT 138.005 82.705 139.215 83.455 ;
        RECT 50.520 82.535 139.300 82.705 ;
        RECT 50.605 81.785 51.815 82.535 ;
        RECT 51.985 81.990 57.330 82.535 ;
        RECT 57.505 81.990 62.850 82.535 ;
        RECT 63.025 81.990 68.370 82.535 ;
        RECT 68.545 81.990 73.890 82.535 ;
        RECT 50.605 81.245 51.125 81.785 ;
        RECT 51.295 81.075 51.815 81.615 ;
        RECT 53.570 81.160 53.910 81.990 ;
        RECT 50.605 79.985 51.815 81.075 ;
        RECT 55.390 80.420 55.740 81.670 ;
        RECT 59.090 81.160 59.430 81.990 ;
        RECT 60.910 80.420 61.260 81.670 ;
        RECT 64.610 81.160 64.950 81.990 ;
        RECT 66.430 80.420 66.780 81.670 ;
        RECT 70.130 81.160 70.470 81.990 ;
        RECT 74.065 81.765 75.735 82.535 ;
        RECT 76.365 81.810 76.655 82.535 ;
        RECT 76.825 81.990 82.170 82.535 ;
        RECT 82.345 81.990 87.690 82.535 ;
        RECT 87.865 81.990 93.210 82.535 ;
        RECT 93.385 81.990 98.730 82.535 ;
        RECT 71.950 80.420 72.300 81.670 ;
        RECT 74.065 81.245 74.815 81.765 ;
        RECT 74.985 81.075 75.735 81.595 ;
        RECT 78.410 81.160 78.750 81.990 ;
        RECT 51.985 79.985 57.330 80.420 ;
        RECT 57.505 79.985 62.850 80.420 ;
        RECT 63.025 79.985 68.370 80.420 ;
        RECT 68.545 79.985 73.890 80.420 ;
        RECT 74.065 79.985 75.735 81.075 ;
        RECT 76.365 79.985 76.655 81.150 ;
        RECT 80.230 80.420 80.580 81.670 ;
        RECT 83.930 81.160 84.270 81.990 ;
        RECT 85.750 80.420 86.100 81.670 ;
        RECT 89.450 81.160 89.790 81.990 ;
        RECT 91.270 80.420 91.620 81.670 ;
        RECT 94.970 81.160 95.310 81.990 ;
        RECT 98.905 81.765 101.495 82.535 ;
        RECT 102.125 81.810 102.415 82.535 ;
        RECT 102.585 81.990 107.930 82.535 ;
        RECT 108.105 81.990 113.450 82.535 ;
        RECT 113.625 81.990 118.970 82.535 ;
        RECT 119.145 81.990 124.490 82.535 ;
        RECT 96.790 80.420 97.140 81.670 ;
        RECT 98.905 81.245 100.115 81.765 ;
        RECT 100.285 81.075 101.495 81.595 ;
        RECT 104.170 81.160 104.510 81.990 ;
        RECT 76.825 79.985 82.170 80.420 ;
        RECT 82.345 79.985 87.690 80.420 ;
        RECT 87.865 79.985 93.210 80.420 ;
        RECT 93.385 79.985 98.730 80.420 ;
        RECT 98.905 79.985 101.495 81.075 ;
        RECT 102.125 79.985 102.415 81.150 ;
        RECT 105.990 80.420 106.340 81.670 ;
        RECT 109.690 81.160 110.030 81.990 ;
        RECT 111.510 80.420 111.860 81.670 ;
        RECT 115.210 81.160 115.550 81.990 ;
        RECT 117.030 80.420 117.380 81.670 ;
        RECT 120.730 81.160 121.070 81.990 ;
        RECT 124.665 81.765 127.255 82.535 ;
        RECT 127.885 81.810 128.175 82.535 ;
        RECT 128.345 81.990 133.690 82.535 ;
        RECT 122.550 80.420 122.900 81.670 ;
        RECT 124.665 81.245 125.875 81.765 ;
        RECT 126.045 81.075 127.255 81.595 ;
        RECT 129.930 81.160 130.270 81.990 ;
        RECT 133.865 81.765 137.375 82.535 ;
        RECT 138.005 81.785 139.215 82.535 ;
        RECT 102.585 79.985 107.930 80.420 ;
        RECT 108.105 79.985 113.450 80.420 ;
        RECT 113.625 79.985 118.970 80.420 ;
        RECT 119.145 79.985 124.490 80.420 ;
        RECT 124.665 79.985 127.255 81.075 ;
        RECT 127.885 79.985 128.175 81.150 ;
        RECT 131.750 80.420 132.100 81.670 ;
        RECT 133.865 81.245 135.515 81.765 ;
        RECT 135.685 81.075 137.375 81.595 ;
        RECT 128.345 79.985 133.690 80.420 ;
        RECT 133.865 79.985 137.375 81.075 ;
        RECT 138.005 81.075 138.525 81.615 ;
        RECT 138.695 81.245 139.215 81.785 ;
        RECT 138.005 79.985 139.215 81.075 ;
        RECT 50.520 79.815 139.300 79.985 ;
        RECT 50.605 78.725 51.815 79.815 ;
        RECT 51.985 79.380 57.330 79.815 ;
        RECT 57.505 79.380 62.850 79.815 ;
        RECT 50.605 78.015 51.125 78.555 ;
        RECT 51.295 78.185 51.815 78.725 ;
        RECT 50.605 77.265 51.815 78.015 ;
        RECT 53.570 77.810 53.910 78.640 ;
        RECT 55.390 78.130 55.740 79.380 ;
        RECT 59.090 77.810 59.430 78.640 ;
        RECT 60.910 78.130 61.260 79.380 ;
        RECT 63.485 78.650 63.775 79.815 ;
        RECT 63.945 79.380 69.290 79.815 ;
        RECT 69.465 79.380 74.810 79.815 ;
        RECT 74.985 79.380 80.330 79.815 ;
        RECT 80.505 79.380 85.850 79.815 ;
        RECT 51.985 77.265 57.330 77.810 ;
        RECT 57.505 77.265 62.850 77.810 ;
        RECT 63.485 77.265 63.775 77.990 ;
        RECT 65.530 77.810 65.870 78.640 ;
        RECT 67.350 78.130 67.700 79.380 ;
        RECT 71.050 77.810 71.390 78.640 ;
        RECT 72.870 78.130 73.220 79.380 ;
        RECT 76.570 77.810 76.910 78.640 ;
        RECT 78.390 78.130 78.740 79.380 ;
        RECT 82.090 77.810 82.430 78.640 ;
        RECT 83.910 78.130 84.260 79.380 ;
        RECT 86.025 78.725 88.615 79.815 ;
        RECT 86.025 78.035 87.235 78.555 ;
        RECT 87.405 78.205 88.615 78.725 ;
        RECT 89.245 78.650 89.535 79.815 ;
        RECT 89.705 79.380 95.050 79.815 ;
        RECT 95.225 79.380 100.570 79.815 ;
        RECT 100.745 79.380 106.090 79.815 ;
        RECT 106.265 79.380 111.610 79.815 ;
        RECT 63.945 77.265 69.290 77.810 ;
        RECT 69.465 77.265 74.810 77.810 ;
        RECT 74.985 77.265 80.330 77.810 ;
        RECT 80.505 77.265 85.850 77.810 ;
        RECT 86.025 77.265 88.615 78.035 ;
        RECT 89.245 77.265 89.535 77.990 ;
        RECT 91.290 77.810 91.630 78.640 ;
        RECT 93.110 78.130 93.460 79.380 ;
        RECT 96.810 77.810 97.150 78.640 ;
        RECT 98.630 78.130 98.980 79.380 ;
        RECT 102.330 77.810 102.670 78.640 ;
        RECT 104.150 78.130 104.500 79.380 ;
        RECT 107.850 77.810 108.190 78.640 ;
        RECT 109.670 78.130 110.020 79.380 ;
        RECT 111.785 78.725 114.375 79.815 ;
        RECT 111.785 78.035 112.995 78.555 ;
        RECT 113.165 78.205 114.375 78.725 ;
        RECT 115.005 78.650 115.295 79.815 ;
        RECT 115.465 79.380 120.810 79.815 ;
        RECT 120.985 79.380 126.330 79.815 ;
        RECT 126.505 79.380 131.850 79.815 ;
        RECT 132.025 79.380 137.370 79.815 ;
        RECT 89.705 77.265 95.050 77.810 ;
        RECT 95.225 77.265 100.570 77.810 ;
        RECT 100.745 77.265 106.090 77.810 ;
        RECT 106.265 77.265 111.610 77.810 ;
        RECT 111.785 77.265 114.375 78.035 ;
        RECT 115.005 77.265 115.295 77.990 ;
        RECT 117.050 77.810 117.390 78.640 ;
        RECT 118.870 78.130 119.220 79.380 ;
        RECT 122.570 77.810 122.910 78.640 ;
        RECT 124.390 78.130 124.740 79.380 ;
        RECT 128.090 77.810 128.430 78.640 ;
        RECT 129.910 78.130 130.260 79.380 ;
        RECT 133.610 77.810 133.950 78.640 ;
        RECT 135.430 78.130 135.780 79.380 ;
        RECT 138.005 78.725 139.215 79.815 ;
        RECT 138.005 78.185 138.525 78.725 ;
        RECT 138.695 78.015 139.215 78.555 ;
        RECT 115.465 77.265 120.810 77.810 ;
        RECT 120.985 77.265 126.330 77.810 ;
        RECT 126.505 77.265 131.850 77.810 ;
        RECT 132.025 77.265 137.370 77.810 ;
        RECT 138.005 77.265 139.215 78.015 ;
        RECT 50.520 77.095 139.300 77.265 ;
        RECT 50.605 76.345 51.815 77.095 ;
        RECT 51.985 76.550 57.330 77.095 ;
        RECT 57.505 76.550 62.850 77.095 ;
        RECT 63.025 76.550 68.370 77.095 ;
        RECT 68.545 76.550 73.890 77.095 ;
        RECT 50.605 75.805 51.125 76.345 ;
        RECT 51.295 75.635 51.815 76.175 ;
        RECT 53.570 75.720 53.910 76.550 ;
        RECT 50.605 74.545 51.815 75.635 ;
        RECT 55.390 74.980 55.740 76.230 ;
        RECT 59.090 75.720 59.430 76.550 ;
        RECT 60.910 74.980 61.260 76.230 ;
        RECT 64.610 75.720 64.950 76.550 ;
        RECT 66.430 74.980 66.780 76.230 ;
        RECT 70.130 75.720 70.470 76.550 ;
        RECT 74.065 76.325 75.735 77.095 ;
        RECT 76.365 76.370 76.655 77.095 ;
        RECT 76.825 76.550 82.170 77.095 ;
        RECT 82.345 76.550 87.690 77.095 ;
        RECT 87.865 76.550 93.210 77.095 ;
        RECT 93.385 76.550 98.730 77.095 ;
        RECT 71.950 74.980 72.300 76.230 ;
        RECT 74.065 75.805 74.815 76.325 ;
        RECT 74.985 75.635 75.735 76.155 ;
        RECT 78.410 75.720 78.750 76.550 ;
        RECT 51.985 74.545 57.330 74.980 ;
        RECT 57.505 74.545 62.850 74.980 ;
        RECT 63.025 74.545 68.370 74.980 ;
        RECT 68.545 74.545 73.890 74.980 ;
        RECT 74.065 74.545 75.735 75.635 ;
        RECT 76.365 74.545 76.655 75.710 ;
        RECT 80.230 74.980 80.580 76.230 ;
        RECT 83.930 75.720 84.270 76.550 ;
        RECT 85.750 74.980 86.100 76.230 ;
        RECT 89.450 75.720 89.790 76.550 ;
        RECT 91.270 74.980 91.620 76.230 ;
        RECT 94.970 75.720 95.310 76.550 ;
        RECT 98.905 76.325 101.495 77.095 ;
        RECT 102.125 76.370 102.415 77.095 ;
        RECT 102.585 76.550 107.930 77.095 ;
        RECT 108.105 76.550 113.450 77.095 ;
        RECT 113.625 76.550 118.970 77.095 ;
        RECT 119.145 76.550 124.490 77.095 ;
        RECT 96.790 74.980 97.140 76.230 ;
        RECT 98.905 75.805 100.115 76.325 ;
        RECT 100.285 75.635 101.495 76.155 ;
        RECT 104.170 75.720 104.510 76.550 ;
        RECT 76.825 74.545 82.170 74.980 ;
        RECT 82.345 74.545 87.690 74.980 ;
        RECT 87.865 74.545 93.210 74.980 ;
        RECT 93.385 74.545 98.730 74.980 ;
        RECT 98.905 74.545 101.495 75.635 ;
        RECT 102.125 74.545 102.415 75.710 ;
        RECT 105.990 74.980 106.340 76.230 ;
        RECT 109.690 75.720 110.030 76.550 ;
        RECT 111.510 74.980 111.860 76.230 ;
        RECT 115.210 75.720 115.550 76.550 ;
        RECT 117.030 74.980 117.380 76.230 ;
        RECT 120.730 75.720 121.070 76.550 ;
        RECT 124.665 76.325 127.255 77.095 ;
        RECT 127.885 76.370 128.175 77.095 ;
        RECT 128.345 76.550 133.690 77.095 ;
        RECT 122.550 74.980 122.900 76.230 ;
        RECT 124.665 75.805 125.875 76.325 ;
        RECT 126.045 75.635 127.255 76.155 ;
        RECT 129.930 75.720 130.270 76.550 ;
        RECT 133.865 76.325 137.375 77.095 ;
        RECT 138.005 76.345 139.215 77.095 ;
        RECT 102.585 74.545 107.930 74.980 ;
        RECT 108.105 74.545 113.450 74.980 ;
        RECT 113.625 74.545 118.970 74.980 ;
        RECT 119.145 74.545 124.490 74.980 ;
        RECT 124.665 74.545 127.255 75.635 ;
        RECT 127.885 74.545 128.175 75.710 ;
        RECT 131.750 74.980 132.100 76.230 ;
        RECT 133.865 75.805 135.515 76.325 ;
        RECT 135.685 75.635 137.375 76.155 ;
        RECT 128.345 74.545 133.690 74.980 ;
        RECT 133.865 74.545 137.375 75.635 ;
        RECT 138.005 75.635 138.525 76.175 ;
        RECT 138.695 75.805 139.215 76.345 ;
        RECT 138.005 74.545 139.215 75.635 ;
        RECT 50.520 74.375 139.300 74.545 ;
        RECT 50.605 73.285 51.815 74.375 ;
        RECT 51.985 73.940 57.330 74.375 ;
        RECT 57.505 73.940 62.850 74.375 ;
        RECT 50.605 72.575 51.125 73.115 ;
        RECT 51.295 72.745 51.815 73.285 ;
        RECT 50.605 71.825 51.815 72.575 ;
        RECT 53.570 72.370 53.910 73.200 ;
        RECT 55.390 72.690 55.740 73.940 ;
        RECT 59.090 72.370 59.430 73.200 ;
        RECT 60.910 72.690 61.260 73.940 ;
        RECT 63.485 73.210 63.775 74.375 ;
        RECT 63.945 73.940 69.290 74.375 ;
        RECT 69.465 73.940 74.810 74.375 ;
        RECT 74.985 73.940 80.330 74.375 ;
        RECT 80.505 73.940 85.850 74.375 ;
        RECT 51.985 71.825 57.330 72.370 ;
        RECT 57.505 71.825 62.850 72.370 ;
        RECT 63.485 71.825 63.775 72.550 ;
        RECT 65.530 72.370 65.870 73.200 ;
        RECT 67.350 72.690 67.700 73.940 ;
        RECT 71.050 72.370 71.390 73.200 ;
        RECT 72.870 72.690 73.220 73.940 ;
        RECT 76.570 72.370 76.910 73.200 ;
        RECT 78.390 72.690 78.740 73.940 ;
        RECT 82.090 72.370 82.430 73.200 ;
        RECT 83.910 72.690 84.260 73.940 ;
        RECT 86.025 73.285 88.615 74.375 ;
        RECT 86.025 72.595 87.235 73.115 ;
        RECT 87.405 72.765 88.615 73.285 ;
        RECT 89.245 73.210 89.535 74.375 ;
        RECT 89.705 73.940 95.050 74.375 ;
        RECT 95.225 73.940 100.570 74.375 ;
        RECT 100.745 73.940 106.090 74.375 ;
        RECT 106.265 73.940 111.610 74.375 ;
        RECT 63.945 71.825 69.290 72.370 ;
        RECT 69.465 71.825 74.810 72.370 ;
        RECT 74.985 71.825 80.330 72.370 ;
        RECT 80.505 71.825 85.850 72.370 ;
        RECT 86.025 71.825 88.615 72.595 ;
        RECT 89.245 71.825 89.535 72.550 ;
        RECT 91.290 72.370 91.630 73.200 ;
        RECT 93.110 72.690 93.460 73.940 ;
        RECT 96.810 72.370 97.150 73.200 ;
        RECT 98.630 72.690 98.980 73.940 ;
        RECT 102.330 72.370 102.670 73.200 ;
        RECT 104.150 72.690 104.500 73.940 ;
        RECT 107.850 72.370 108.190 73.200 ;
        RECT 109.670 72.690 110.020 73.940 ;
        RECT 111.785 73.285 114.375 74.375 ;
        RECT 111.785 72.595 112.995 73.115 ;
        RECT 113.165 72.765 114.375 73.285 ;
        RECT 115.005 73.210 115.295 74.375 ;
        RECT 115.465 73.940 120.810 74.375 ;
        RECT 120.985 73.940 126.330 74.375 ;
        RECT 126.505 73.940 131.850 74.375 ;
        RECT 132.025 73.940 137.370 74.375 ;
        RECT 89.705 71.825 95.050 72.370 ;
        RECT 95.225 71.825 100.570 72.370 ;
        RECT 100.745 71.825 106.090 72.370 ;
        RECT 106.265 71.825 111.610 72.370 ;
        RECT 111.785 71.825 114.375 72.595 ;
        RECT 115.005 71.825 115.295 72.550 ;
        RECT 117.050 72.370 117.390 73.200 ;
        RECT 118.870 72.690 119.220 73.940 ;
        RECT 122.570 72.370 122.910 73.200 ;
        RECT 124.390 72.690 124.740 73.940 ;
        RECT 128.090 72.370 128.430 73.200 ;
        RECT 129.910 72.690 130.260 73.940 ;
        RECT 133.610 72.370 133.950 73.200 ;
        RECT 135.430 72.690 135.780 73.940 ;
        RECT 138.005 73.285 139.215 74.375 ;
        RECT 138.005 72.745 138.525 73.285 ;
        RECT 138.695 72.575 139.215 73.115 ;
        RECT 115.465 71.825 120.810 72.370 ;
        RECT 120.985 71.825 126.330 72.370 ;
        RECT 126.505 71.825 131.850 72.370 ;
        RECT 132.025 71.825 137.370 72.370 ;
        RECT 138.005 71.825 139.215 72.575 ;
        RECT 50.520 71.655 139.300 71.825 ;
        RECT 50.605 70.905 51.815 71.655 ;
        RECT 51.985 71.110 57.330 71.655 ;
        RECT 57.505 71.110 62.850 71.655 ;
        RECT 63.025 71.110 68.370 71.655 ;
        RECT 68.545 71.110 73.890 71.655 ;
        RECT 50.605 70.365 51.125 70.905 ;
        RECT 51.295 70.195 51.815 70.735 ;
        RECT 53.570 70.280 53.910 71.110 ;
        RECT 50.605 69.105 51.815 70.195 ;
        RECT 55.390 69.540 55.740 70.790 ;
        RECT 59.090 70.280 59.430 71.110 ;
        RECT 60.910 69.540 61.260 70.790 ;
        RECT 64.610 70.280 64.950 71.110 ;
        RECT 66.430 69.540 66.780 70.790 ;
        RECT 70.130 70.280 70.470 71.110 ;
        RECT 74.065 70.885 75.735 71.655 ;
        RECT 76.365 70.930 76.655 71.655 ;
        RECT 76.825 71.110 82.170 71.655 ;
        RECT 82.345 71.110 87.690 71.655 ;
        RECT 87.865 71.110 93.210 71.655 ;
        RECT 93.385 71.110 98.730 71.655 ;
        RECT 71.950 69.540 72.300 70.790 ;
        RECT 74.065 70.365 74.815 70.885 ;
        RECT 74.985 70.195 75.735 70.715 ;
        RECT 78.410 70.280 78.750 71.110 ;
        RECT 51.985 69.105 57.330 69.540 ;
        RECT 57.505 69.105 62.850 69.540 ;
        RECT 63.025 69.105 68.370 69.540 ;
        RECT 68.545 69.105 73.890 69.540 ;
        RECT 74.065 69.105 75.735 70.195 ;
        RECT 76.365 69.105 76.655 70.270 ;
        RECT 80.230 69.540 80.580 70.790 ;
        RECT 83.930 70.280 84.270 71.110 ;
        RECT 85.750 69.540 86.100 70.790 ;
        RECT 89.450 70.280 89.790 71.110 ;
        RECT 91.270 69.540 91.620 70.790 ;
        RECT 94.970 70.280 95.310 71.110 ;
        RECT 98.905 70.885 101.495 71.655 ;
        RECT 102.125 70.930 102.415 71.655 ;
        RECT 102.585 71.110 107.930 71.655 ;
        RECT 108.105 71.110 113.450 71.655 ;
        RECT 113.625 71.110 118.970 71.655 ;
        RECT 119.145 71.110 124.490 71.655 ;
        RECT 96.790 69.540 97.140 70.790 ;
        RECT 98.905 70.365 100.115 70.885 ;
        RECT 100.285 70.195 101.495 70.715 ;
        RECT 104.170 70.280 104.510 71.110 ;
        RECT 76.825 69.105 82.170 69.540 ;
        RECT 82.345 69.105 87.690 69.540 ;
        RECT 87.865 69.105 93.210 69.540 ;
        RECT 93.385 69.105 98.730 69.540 ;
        RECT 98.905 69.105 101.495 70.195 ;
        RECT 102.125 69.105 102.415 70.270 ;
        RECT 105.990 69.540 106.340 70.790 ;
        RECT 109.690 70.280 110.030 71.110 ;
        RECT 111.510 69.540 111.860 70.790 ;
        RECT 115.210 70.280 115.550 71.110 ;
        RECT 117.030 69.540 117.380 70.790 ;
        RECT 120.730 70.280 121.070 71.110 ;
        RECT 124.665 70.885 127.255 71.655 ;
        RECT 127.885 70.930 128.175 71.655 ;
        RECT 128.345 71.110 133.690 71.655 ;
        RECT 122.550 69.540 122.900 70.790 ;
        RECT 124.665 70.365 125.875 70.885 ;
        RECT 126.045 70.195 127.255 70.715 ;
        RECT 129.930 70.280 130.270 71.110 ;
        RECT 133.865 70.885 137.375 71.655 ;
        RECT 138.005 70.905 139.215 71.655 ;
        RECT 102.585 69.105 107.930 69.540 ;
        RECT 108.105 69.105 113.450 69.540 ;
        RECT 113.625 69.105 118.970 69.540 ;
        RECT 119.145 69.105 124.490 69.540 ;
        RECT 124.665 69.105 127.255 70.195 ;
        RECT 127.885 69.105 128.175 70.270 ;
        RECT 131.750 69.540 132.100 70.790 ;
        RECT 133.865 70.365 135.515 70.885 ;
        RECT 135.685 70.195 137.375 70.715 ;
        RECT 128.345 69.105 133.690 69.540 ;
        RECT 133.865 69.105 137.375 70.195 ;
        RECT 138.005 70.195 138.525 70.735 ;
        RECT 138.695 70.365 139.215 70.905 ;
        RECT 138.005 69.105 139.215 70.195 ;
        RECT 50.520 68.935 139.300 69.105 ;
        RECT 50.605 67.845 51.815 68.935 ;
        RECT 51.985 68.500 57.330 68.935 ;
        RECT 57.505 68.500 62.850 68.935 ;
        RECT 50.605 67.135 51.125 67.675 ;
        RECT 51.295 67.305 51.815 67.845 ;
        RECT 50.605 66.385 51.815 67.135 ;
        RECT 53.570 66.930 53.910 67.760 ;
        RECT 55.390 67.250 55.740 68.500 ;
        RECT 59.090 66.930 59.430 67.760 ;
        RECT 60.910 67.250 61.260 68.500 ;
        RECT 63.485 67.770 63.775 68.935 ;
        RECT 63.945 68.500 69.290 68.935 ;
        RECT 69.465 68.500 74.810 68.935 ;
        RECT 74.985 68.500 80.330 68.935 ;
        RECT 80.505 68.500 85.850 68.935 ;
        RECT 51.985 66.385 57.330 66.930 ;
        RECT 57.505 66.385 62.850 66.930 ;
        RECT 63.485 66.385 63.775 67.110 ;
        RECT 65.530 66.930 65.870 67.760 ;
        RECT 67.350 67.250 67.700 68.500 ;
        RECT 71.050 66.930 71.390 67.760 ;
        RECT 72.870 67.250 73.220 68.500 ;
        RECT 76.570 66.930 76.910 67.760 ;
        RECT 78.390 67.250 78.740 68.500 ;
        RECT 82.090 66.930 82.430 67.760 ;
        RECT 83.910 67.250 84.260 68.500 ;
        RECT 86.025 67.845 88.615 68.935 ;
        RECT 86.025 67.155 87.235 67.675 ;
        RECT 87.405 67.325 88.615 67.845 ;
        RECT 89.245 67.770 89.535 68.935 ;
        RECT 89.705 68.500 95.050 68.935 ;
        RECT 95.225 68.500 100.570 68.935 ;
        RECT 100.745 68.500 106.090 68.935 ;
        RECT 106.265 68.500 111.610 68.935 ;
        RECT 63.945 66.385 69.290 66.930 ;
        RECT 69.465 66.385 74.810 66.930 ;
        RECT 74.985 66.385 80.330 66.930 ;
        RECT 80.505 66.385 85.850 66.930 ;
        RECT 86.025 66.385 88.615 67.155 ;
        RECT 89.245 66.385 89.535 67.110 ;
        RECT 91.290 66.930 91.630 67.760 ;
        RECT 93.110 67.250 93.460 68.500 ;
        RECT 96.810 66.930 97.150 67.760 ;
        RECT 98.630 67.250 98.980 68.500 ;
        RECT 102.330 66.930 102.670 67.760 ;
        RECT 104.150 67.250 104.500 68.500 ;
        RECT 107.850 66.930 108.190 67.760 ;
        RECT 109.670 67.250 110.020 68.500 ;
        RECT 111.785 67.845 114.375 68.935 ;
        RECT 111.785 67.155 112.995 67.675 ;
        RECT 113.165 67.325 114.375 67.845 ;
        RECT 115.005 67.770 115.295 68.935 ;
        RECT 115.465 68.500 120.810 68.935 ;
        RECT 120.985 68.500 126.330 68.935 ;
        RECT 126.505 68.500 131.850 68.935 ;
        RECT 132.025 68.500 137.370 68.935 ;
        RECT 89.705 66.385 95.050 66.930 ;
        RECT 95.225 66.385 100.570 66.930 ;
        RECT 100.745 66.385 106.090 66.930 ;
        RECT 106.265 66.385 111.610 66.930 ;
        RECT 111.785 66.385 114.375 67.155 ;
        RECT 115.005 66.385 115.295 67.110 ;
        RECT 117.050 66.930 117.390 67.760 ;
        RECT 118.870 67.250 119.220 68.500 ;
        RECT 122.570 66.930 122.910 67.760 ;
        RECT 124.390 67.250 124.740 68.500 ;
        RECT 128.090 66.930 128.430 67.760 ;
        RECT 129.910 67.250 130.260 68.500 ;
        RECT 133.610 66.930 133.950 67.760 ;
        RECT 135.430 67.250 135.780 68.500 ;
        RECT 138.005 67.845 139.215 68.935 ;
        RECT 138.005 67.305 138.525 67.845 ;
        RECT 138.695 67.135 139.215 67.675 ;
        RECT 115.465 66.385 120.810 66.930 ;
        RECT 120.985 66.385 126.330 66.930 ;
        RECT 126.505 66.385 131.850 66.930 ;
        RECT 132.025 66.385 137.370 66.930 ;
        RECT 138.005 66.385 139.215 67.135 ;
        RECT 50.520 66.215 139.300 66.385 ;
        RECT 50.605 65.465 51.815 66.215 ;
        RECT 51.985 65.670 57.330 66.215 ;
        RECT 57.505 65.670 62.850 66.215 ;
        RECT 63.025 65.670 68.370 66.215 ;
        RECT 68.545 65.670 73.890 66.215 ;
        RECT 50.605 64.925 51.125 65.465 ;
        RECT 51.295 64.755 51.815 65.295 ;
        RECT 53.570 64.840 53.910 65.670 ;
        RECT 50.605 63.665 51.815 64.755 ;
        RECT 55.390 64.100 55.740 65.350 ;
        RECT 59.090 64.840 59.430 65.670 ;
        RECT 60.910 64.100 61.260 65.350 ;
        RECT 64.610 64.840 64.950 65.670 ;
        RECT 66.430 64.100 66.780 65.350 ;
        RECT 70.130 64.840 70.470 65.670 ;
        RECT 74.065 65.445 75.735 66.215 ;
        RECT 76.365 65.490 76.655 66.215 ;
        RECT 76.825 65.670 82.170 66.215 ;
        RECT 82.345 65.670 87.690 66.215 ;
        RECT 87.865 65.670 93.210 66.215 ;
        RECT 93.385 65.670 98.730 66.215 ;
        RECT 71.950 64.100 72.300 65.350 ;
        RECT 74.065 64.925 74.815 65.445 ;
        RECT 74.985 64.755 75.735 65.275 ;
        RECT 78.410 64.840 78.750 65.670 ;
        RECT 51.985 63.665 57.330 64.100 ;
        RECT 57.505 63.665 62.850 64.100 ;
        RECT 63.025 63.665 68.370 64.100 ;
        RECT 68.545 63.665 73.890 64.100 ;
        RECT 74.065 63.665 75.735 64.755 ;
        RECT 76.365 63.665 76.655 64.830 ;
        RECT 80.230 64.100 80.580 65.350 ;
        RECT 83.930 64.840 84.270 65.670 ;
        RECT 85.750 64.100 86.100 65.350 ;
        RECT 89.450 64.840 89.790 65.670 ;
        RECT 91.270 64.100 91.620 65.350 ;
        RECT 94.970 64.840 95.310 65.670 ;
        RECT 98.905 65.445 101.495 66.215 ;
        RECT 102.125 65.490 102.415 66.215 ;
        RECT 102.585 65.670 107.930 66.215 ;
        RECT 108.105 65.670 113.450 66.215 ;
        RECT 113.625 65.670 118.970 66.215 ;
        RECT 119.145 65.670 124.490 66.215 ;
        RECT 96.790 64.100 97.140 65.350 ;
        RECT 98.905 64.925 100.115 65.445 ;
        RECT 100.285 64.755 101.495 65.275 ;
        RECT 104.170 64.840 104.510 65.670 ;
        RECT 76.825 63.665 82.170 64.100 ;
        RECT 82.345 63.665 87.690 64.100 ;
        RECT 87.865 63.665 93.210 64.100 ;
        RECT 93.385 63.665 98.730 64.100 ;
        RECT 98.905 63.665 101.495 64.755 ;
        RECT 102.125 63.665 102.415 64.830 ;
        RECT 105.990 64.100 106.340 65.350 ;
        RECT 109.690 64.840 110.030 65.670 ;
        RECT 111.510 64.100 111.860 65.350 ;
        RECT 115.210 64.840 115.550 65.670 ;
        RECT 117.030 64.100 117.380 65.350 ;
        RECT 120.730 64.840 121.070 65.670 ;
        RECT 124.665 65.445 127.255 66.215 ;
        RECT 127.885 65.490 128.175 66.215 ;
        RECT 128.345 65.670 133.690 66.215 ;
        RECT 122.550 64.100 122.900 65.350 ;
        RECT 124.665 64.925 125.875 65.445 ;
        RECT 126.045 64.755 127.255 65.275 ;
        RECT 129.930 64.840 130.270 65.670 ;
        RECT 133.865 65.445 137.375 66.215 ;
        RECT 138.005 65.465 139.215 66.215 ;
        RECT 102.585 63.665 107.930 64.100 ;
        RECT 108.105 63.665 113.450 64.100 ;
        RECT 113.625 63.665 118.970 64.100 ;
        RECT 119.145 63.665 124.490 64.100 ;
        RECT 124.665 63.665 127.255 64.755 ;
        RECT 127.885 63.665 128.175 64.830 ;
        RECT 131.750 64.100 132.100 65.350 ;
        RECT 133.865 64.925 135.515 65.445 ;
        RECT 135.685 64.755 137.375 65.275 ;
        RECT 128.345 63.665 133.690 64.100 ;
        RECT 133.865 63.665 137.375 64.755 ;
        RECT 138.005 64.755 138.525 65.295 ;
        RECT 138.695 64.925 139.215 65.465 ;
        RECT 138.005 63.665 139.215 64.755 ;
        RECT 50.520 63.495 139.300 63.665 ;
        RECT 50.605 62.405 51.815 63.495 ;
        RECT 51.985 63.060 57.330 63.495 ;
        RECT 57.505 63.060 62.850 63.495 ;
        RECT 50.605 61.695 51.125 62.235 ;
        RECT 51.295 61.865 51.815 62.405 ;
        RECT 50.605 60.945 51.815 61.695 ;
        RECT 53.570 61.490 53.910 62.320 ;
        RECT 55.390 61.810 55.740 63.060 ;
        RECT 59.090 61.490 59.430 62.320 ;
        RECT 60.910 61.810 61.260 63.060 ;
        RECT 63.485 62.330 63.775 63.495 ;
        RECT 63.945 63.060 69.290 63.495 ;
        RECT 69.465 63.060 74.810 63.495 ;
        RECT 51.985 60.945 57.330 61.490 ;
        RECT 57.505 60.945 62.850 61.490 ;
        RECT 63.485 60.945 63.775 61.670 ;
        RECT 65.530 61.490 65.870 62.320 ;
        RECT 67.350 61.810 67.700 63.060 ;
        RECT 71.050 61.490 71.390 62.320 ;
        RECT 72.870 61.810 73.220 63.060 ;
        RECT 74.985 62.405 76.195 63.495 ;
        RECT 74.985 61.695 75.505 62.235 ;
        RECT 75.675 61.865 76.195 62.405 ;
        RECT 76.365 62.330 76.655 63.495 ;
        RECT 76.825 63.060 82.170 63.495 ;
        RECT 82.345 63.060 87.690 63.495 ;
        RECT 63.945 60.945 69.290 61.490 ;
        RECT 69.465 60.945 74.810 61.490 ;
        RECT 74.985 60.945 76.195 61.695 ;
        RECT 76.365 60.945 76.655 61.670 ;
        RECT 78.410 61.490 78.750 62.320 ;
        RECT 80.230 61.810 80.580 63.060 ;
        RECT 83.930 61.490 84.270 62.320 ;
        RECT 85.750 61.810 86.100 63.060 ;
        RECT 87.865 62.405 89.075 63.495 ;
        RECT 87.865 61.695 88.385 62.235 ;
        RECT 88.555 61.865 89.075 62.405 ;
        RECT 89.245 62.330 89.535 63.495 ;
        RECT 89.705 63.060 95.050 63.495 ;
        RECT 95.225 63.060 100.570 63.495 ;
        RECT 76.825 60.945 82.170 61.490 ;
        RECT 82.345 60.945 87.690 61.490 ;
        RECT 87.865 60.945 89.075 61.695 ;
        RECT 89.245 60.945 89.535 61.670 ;
        RECT 91.290 61.490 91.630 62.320 ;
        RECT 93.110 61.810 93.460 63.060 ;
        RECT 96.810 61.490 97.150 62.320 ;
        RECT 98.630 61.810 98.980 63.060 ;
        RECT 100.745 62.405 101.955 63.495 ;
        RECT 100.745 61.695 101.265 62.235 ;
        RECT 101.435 61.865 101.955 62.405 ;
        RECT 102.125 62.330 102.415 63.495 ;
        RECT 102.585 63.060 107.930 63.495 ;
        RECT 108.105 63.060 113.450 63.495 ;
        RECT 89.705 60.945 95.050 61.490 ;
        RECT 95.225 60.945 100.570 61.490 ;
        RECT 100.745 60.945 101.955 61.695 ;
        RECT 102.125 60.945 102.415 61.670 ;
        RECT 104.170 61.490 104.510 62.320 ;
        RECT 105.990 61.810 106.340 63.060 ;
        RECT 109.690 61.490 110.030 62.320 ;
        RECT 111.510 61.810 111.860 63.060 ;
        RECT 113.625 62.405 114.835 63.495 ;
        RECT 113.625 61.695 114.145 62.235 ;
        RECT 114.315 61.865 114.835 62.405 ;
        RECT 115.005 62.330 115.295 63.495 ;
        RECT 115.465 63.060 120.810 63.495 ;
        RECT 120.985 63.060 126.330 63.495 ;
        RECT 102.585 60.945 107.930 61.490 ;
        RECT 108.105 60.945 113.450 61.490 ;
        RECT 113.625 60.945 114.835 61.695 ;
        RECT 115.005 60.945 115.295 61.670 ;
        RECT 117.050 61.490 117.390 62.320 ;
        RECT 118.870 61.810 119.220 63.060 ;
        RECT 122.570 61.490 122.910 62.320 ;
        RECT 124.390 61.810 124.740 63.060 ;
        RECT 126.505 62.405 127.715 63.495 ;
        RECT 126.505 61.695 127.025 62.235 ;
        RECT 127.195 61.865 127.715 62.405 ;
        RECT 127.885 62.330 128.175 63.495 ;
        RECT 128.345 63.060 133.690 63.495 ;
        RECT 115.465 60.945 120.810 61.490 ;
        RECT 120.985 60.945 126.330 61.490 ;
        RECT 126.505 60.945 127.715 61.695 ;
        RECT 127.885 60.945 128.175 61.670 ;
        RECT 129.930 61.490 130.270 62.320 ;
        RECT 131.750 61.810 132.100 63.060 ;
        RECT 133.865 62.405 137.375 63.495 ;
        RECT 133.865 61.715 135.515 62.235 ;
        RECT 135.685 61.885 137.375 62.405 ;
        RECT 138.005 62.405 139.215 63.495 ;
        RECT 138.005 61.865 138.525 62.405 ;
        RECT 128.345 60.945 133.690 61.490 ;
        RECT 133.865 60.945 137.375 61.715 ;
        RECT 138.695 61.695 139.215 62.235 ;
        RECT 138.005 60.945 139.215 61.695 ;
        RECT 50.520 60.775 139.300 60.945 ;
      LAYER mcon ;
        RECT 50.665 136.935 50.835 137.105 ;
        RECT 51.125 136.935 51.295 137.105 ;
        RECT 51.585 136.935 51.755 137.105 ;
        RECT 52.045 136.935 52.215 137.105 ;
        RECT 52.505 136.935 52.675 137.105 ;
        RECT 52.965 136.935 53.135 137.105 ;
        RECT 53.425 136.935 53.595 137.105 ;
        RECT 53.885 136.935 54.055 137.105 ;
        RECT 54.345 136.935 54.515 137.105 ;
        RECT 54.805 136.935 54.975 137.105 ;
        RECT 55.265 136.935 55.435 137.105 ;
        RECT 55.725 136.935 55.895 137.105 ;
        RECT 56.185 136.935 56.355 137.105 ;
        RECT 56.645 136.935 56.815 137.105 ;
        RECT 57.105 136.935 57.275 137.105 ;
        RECT 57.565 136.935 57.735 137.105 ;
        RECT 58.025 136.935 58.195 137.105 ;
        RECT 58.485 136.935 58.655 137.105 ;
        RECT 58.945 136.935 59.115 137.105 ;
        RECT 59.405 136.935 59.575 137.105 ;
        RECT 59.865 136.935 60.035 137.105 ;
        RECT 60.325 136.935 60.495 137.105 ;
        RECT 60.785 136.935 60.955 137.105 ;
        RECT 61.245 136.935 61.415 137.105 ;
        RECT 61.705 136.935 61.875 137.105 ;
        RECT 62.165 136.935 62.335 137.105 ;
        RECT 62.625 136.935 62.795 137.105 ;
        RECT 63.085 136.935 63.255 137.105 ;
        RECT 63.545 136.935 63.715 137.105 ;
        RECT 64.005 136.935 64.175 137.105 ;
        RECT 64.465 136.935 64.635 137.105 ;
        RECT 64.925 136.935 65.095 137.105 ;
        RECT 65.385 136.935 65.555 137.105 ;
        RECT 65.845 136.935 66.015 137.105 ;
        RECT 66.305 136.935 66.475 137.105 ;
        RECT 66.765 136.935 66.935 137.105 ;
        RECT 67.225 136.935 67.395 137.105 ;
        RECT 67.685 136.935 67.855 137.105 ;
        RECT 68.145 136.935 68.315 137.105 ;
        RECT 68.605 136.935 68.775 137.105 ;
        RECT 69.065 136.935 69.235 137.105 ;
        RECT 69.525 136.935 69.695 137.105 ;
        RECT 69.985 136.935 70.155 137.105 ;
        RECT 70.445 136.935 70.615 137.105 ;
        RECT 70.905 136.935 71.075 137.105 ;
        RECT 71.365 136.935 71.535 137.105 ;
        RECT 71.825 136.935 71.995 137.105 ;
        RECT 72.285 136.935 72.455 137.105 ;
        RECT 72.745 136.935 72.915 137.105 ;
        RECT 73.205 136.935 73.375 137.105 ;
        RECT 73.665 136.935 73.835 137.105 ;
        RECT 74.125 136.935 74.295 137.105 ;
        RECT 74.585 136.935 74.755 137.105 ;
        RECT 75.045 136.935 75.215 137.105 ;
        RECT 75.505 136.935 75.675 137.105 ;
        RECT 75.965 136.935 76.135 137.105 ;
        RECT 76.425 136.935 76.595 137.105 ;
        RECT 76.885 136.935 77.055 137.105 ;
        RECT 77.345 136.935 77.515 137.105 ;
        RECT 77.805 136.935 77.975 137.105 ;
        RECT 78.265 136.935 78.435 137.105 ;
        RECT 78.725 136.935 78.895 137.105 ;
        RECT 79.185 136.935 79.355 137.105 ;
        RECT 79.645 136.935 79.815 137.105 ;
        RECT 80.105 136.935 80.275 137.105 ;
        RECT 80.565 136.935 80.735 137.105 ;
        RECT 81.025 136.935 81.195 137.105 ;
        RECT 81.485 136.935 81.655 137.105 ;
        RECT 81.945 136.935 82.115 137.105 ;
        RECT 82.405 136.935 82.575 137.105 ;
        RECT 82.865 136.935 83.035 137.105 ;
        RECT 83.325 136.935 83.495 137.105 ;
        RECT 83.785 136.935 83.955 137.105 ;
        RECT 84.245 136.935 84.415 137.105 ;
        RECT 84.705 136.935 84.875 137.105 ;
        RECT 85.165 136.935 85.335 137.105 ;
        RECT 85.625 136.935 85.795 137.105 ;
        RECT 86.085 136.935 86.255 137.105 ;
        RECT 86.545 136.935 86.715 137.105 ;
        RECT 87.005 136.935 87.175 137.105 ;
        RECT 87.465 136.935 87.635 137.105 ;
        RECT 87.925 136.935 88.095 137.105 ;
        RECT 88.385 136.935 88.555 137.105 ;
        RECT 88.845 136.935 89.015 137.105 ;
        RECT 89.305 136.935 89.475 137.105 ;
        RECT 89.765 136.935 89.935 137.105 ;
        RECT 90.225 136.935 90.395 137.105 ;
        RECT 90.685 136.935 90.855 137.105 ;
        RECT 91.145 136.935 91.315 137.105 ;
        RECT 91.605 136.935 91.775 137.105 ;
        RECT 92.065 136.935 92.235 137.105 ;
        RECT 92.525 136.935 92.695 137.105 ;
        RECT 92.985 136.935 93.155 137.105 ;
        RECT 93.445 136.935 93.615 137.105 ;
        RECT 93.905 136.935 94.075 137.105 ;
        RECT 94.365 136.935 94.535 137.105 ;
        RECT 94.825 136.935 94.995 137.105 ;
        RECT 95.285 136.935 95.455 137.105 ;
        RECT 95.745 136.935 95.915 137.105 ;
        RECT 96.205 136.935 96.375 137.105 ;
        RECT 96.665 136.935 96.835 137.105 ;
        RECT 97.125 136.935 97.295 137.105 ;
        RECT 97.585 136.935 97.755 137.105 ;
        RECT 98.045 136.935 98.215 137.105 ;
        RECT 98.505 136.935 98.675 137.105 ;
        RECT 98.965 136.935 99.135 137.105 ;
        RECT 99.425 136.935 99.595 137.105 ;
        RECT 99.885 136.935 100.055 137.105 ;
        RECT 100.345 136.935 100.515 137.105 ;
        RECT 100.805 136.935 100.975 137.105 ;
        RECT 101.265 136.935 101.435 137.105 ;
        RECT 101.725 136.935 101.895 137.105 ;
        RECT 102.185 136.935 102.355 137.105 ;
        RECT 102.645 136.935 102.815 137.105 ;
        RECT 103.105 136.935 103.275 137.105 ;
        RECT 103.565 136.935 103.735 137.105 ;
        RECT 104.025 136.935 104.195 137.105 ;
        RECT 104.485 136.935 104.655 137.105 ;
        RECT 104.945 136.935 105.115 137.105 ;
        RECT 105.405 136.935 105.575 137.105 ;
        RECT 105.865 136.935 106.035 137.105 ;
        RECT 106.325 136.935 106.495 137.105 ;
        RECT 106.785 136.935 106.955 137.105 ;
        RECT 107.245 136.935 107.415 137.105 ;
        RECT 107.705 136.935 107.875 137.105 ;
        RECT 108.165 136.935 108.335 137.105 ;
        RECT 108.625 136.935 108.795 137.105 ;
        RECT 109.085 136.935 109.255 137.105 ;
        RECT 109.545 136.935 109.715 137.105 ;
        RECT 110.005 136.935 110.175 137.105 ;
        RECT 110.465 136.935 110.635 137.105 ;
        RECT 110.925 136.935 111.095 137.105 ;
        RECT 111.385 136.935 111.555 137.105 ;
        RECT 111.845 136.935 112.015 137.105 ;
        RECT 112.305 136.935 112.475 137.105 ;
        RECT 112.765 136.935 112.935 137.105 ;
        RECT 113.225 136.935 113.395 137.105 ;
        RECT 113.685 136.935 113.855 137.105 ;
        RECT 114.145 136.935 114.315 137.105 ;
        RECT 114.605 136.935 114.775 137.105 ;
        RECT 115.065 136.935 115.235 137.105 ;
        RECT 115.525 136.935 115.695 137.105 ;
        RECT 115.985 136.935 116.155 137.105 ;
        RECT 116.445 136.935 116.615 137.105 ;
        RECT 116.905 136.935 117.075 137.105 ;
        RECT 117.365 136.935 117.535 137.105 ;
        RECT 117.825 136.935 117.995 137.105 ;
        RECT 118.285 136.935 118.455 137.105 ;
        RECT 118.745 136.935 118.915 137.105 ;
        RECT 119.205 136.935 119.375 137.105 ;
        RECT 119.665 136.935 119.835 137.105 ;
        RECT 120.125 136.935 120.295 137.105 ;
        RECT 120.585 136.935 120.755 137.105 ;
        RECT 121.045 136.935 121.215 137.105 ;
        RECT 121.505 136.935 121.675 137.105 ;
        RECT 121.965 136.935 122.135 137.105 ;
        RECT 122.425 136.935 122.595 137.105 ;
        RECT 122.885 136.935 123.055 137.105 ;
        RECT 123.345 136.935 123.515 137.105 ;
        RECT 123.805 136.935 123.975 137.105 ;
        RECT 124.265 136.935 124.435 137.105 ;
        RECT 124.725 136.935 124.895 137.105 ;
        RECT 125.185 136.935 125.355 137.105 ;
        RECT 125.645 136.935 125.815 137.105 ;
        RECT 126.105 136.935 126.275 137.105 ;
        RECT 126.565 136.935 126.735 137.105 ;
        RECT 127.025 136.935 127.195 137.105 ;
        RECT 127.485 136.935 127.655 137.105 ;
        RECT 127.945 136.935 128.115 137.105 ;
        RECT 128.405 136.935 128.575 137.105 ;
        RECT 128.865 136.935 129.035 137.105 ;
        RECT 129.325 136.935 129.495 137.105 ;
        RECT 129.785 136.935 129.955 137.105 ;
        RECT 130.245 136.935 130.415 137.105 ;
        RECT 130.705 136.935 130.875 137.105 ;
        RECT 131.165 136.935 131.335 137.105 ;
        RECT 131.625 136.935 131.795 137.105 ;
        RECT 132.085 136.935 132.255 137.105 ;
        RECT 132.545 136.935 132.715 137.105 ;
        RECT 133.005 136.935 133.175 137.105 ;
        RECT 133.465 136.935 133.635 137.105 ;
        RECT 133.925 136.935 134.095 137.105 ;
        RECT 134.385 136.935 134.555 137.105 ;
        RECT 134.845 136.935 135.015 137.105 ;
        RECT 135.305 136.935 135.475 137.105 ;
        RECT 135.765 136.935 135.935 137.105 ;
        RECT 136.225 136.935 136.395 137.105 ;
        RECT 136.685 136.935 136.855 137.105 ;
        RECT 137.145 136.935 137.315 137.105 ;
        RECT 137.605 136.935 137.775 137.105 ;
        RECT 138.065 136.935 138.235 137.105 ;
        RECT 138.525 136.935 138.695 137.105 ;
        RECT 138.985 136.935 139.155 137.105 ;
        RECT 50.665 134.215 50.835 134.385 ;
        RECT 51.125 134.215 51.295 134.385 ;
        RECT 51.585 134.215 51.755 134.385 ;
        RECT 52.045 134.215 52.215 134.385 ;
        RECT 52.505 134.215 52.675 134.385 ;
        RECT 52.965 134.215 53.135 134.385 ;
        RECT 53.425 134.215 53.595 134.385 ;
        RECT 53.885 134.215 54.055 134.385 ;
        RECT 54.345 134.215 54.515 134.385 ;
        RECT 54.805 134.215 54.975 134.385 ;
        RECT 55.265 134.215 55.435 134.385 ;
        RECT 55.725 134.215 55.895 134.385 ;
        RECT 56.185 134.215 56.355 134.385 ;
        RECT 56.645 134.215 56.815 134.385 ;
        RECT 57.105 134.215 57.275 134.385 ;
        RECT 57.565 134.215 57.735 134.385 ;
        RECT 58.025 134.215 58.195 134.385 ;
        RECT 58.485 134.215 58.655 134.385 ;
        RECT 58.945 134.215 59.115 134.385 ;
        RECT 59.405 134.215 59.575 134.385 ;
        RECT 59.865 134.215 60.035 134.385 ;
        RECT 60.325 134.215 60.495 134.385 ;
        RECT 60.785 134.215 60.955 134.385 ;
        RECT 61.245 134.215 61.415 134.385 ;
        RECT 61.705 134.215 61.875 134.385 ;
        RECT 62.165 134.215 62.335 134.385 ;
        RECT 62.625 134.215 62.795 134.385 ;
        RECT 63.085 134.215 63.255 134.385 ;
        RECT 63.545 134.215 63.715 134.385 ;
        RECT 64.005 134.215 64.175 134.385 ;
        RECT 64.465 134.215 64.635 134.385 ;
        RECT 64.925 134.215 65.095 134.385 ;
        RECT 65.385 134.215 65.555 134.385 ;
        RECT 65.845 134.215 66.015 134.385 ;
        RECT 66.305 134.215 66.475 134.385 ;
        RECT 66.765 134.215 66.935 134.385 ;
        RECT 67.225 134.215 67.395 134.385 ;
        RECT 67.685 134.215 67.855 134.385 ;
        RECT 68.145 134.215 68.315 134.385 ;
        RECT 68.605 134.215 68.775 134.385 ;
        RECT 69.065 134.215 69.235 134.385 ;
        RECT 69.525 134.215 69.695 134.385 ;
        RECT 69.985 134.215 70.155 134.385 ;
        RECT 70.445 134.215 70.615 134.385 ;
        RECT 70.905 134.215 71.075 134.385 ;
        RECT 71.365 134.215 71.535 134.385 ;
        RECT 71.825 134.215 71.995 134.385 ;
        RECT 72.285 134.215 72.455 134.385 ;
        RECT 72.745 134.215 72.915 134.385 ;
        RECT 73.205 134.215 73.375 134.385 ;
        RECT 73.665 134.215 73.835 134.385 ;
        RECT 74.125 134.215 74.295 134.385 ;
        RECT 74.585 134.215 74.755 134.385 ;
        RECT 75.045 134.215 75.215 134.385 ;
        RECT 75.505 134.215 75.675 134.385 ;
        RECT 75.965 134.215 76.135 134.385 ;
        RECT 76.425 134.215 76.595 134.385 ;
        RECT 76.885 134.215 77.055 134.385 ;
        RECT 77.345 134.215 77.515 134.385 ;
        RECT 77.805 134.215 77.975 134.385 ;
        RECT 78.265 134.215 78.435 134.385 ;
        RECT 78.725 134.215 78.895 134.385 ;
        RECT 79.185 134.215 79.355 134.385 ;
        RECT 79.645 134.215 79.815 134.385 ;
        RECT 80.105 134.215 80.275 134.385 ;
        RECT 80.565 134.215 80.735 134.385 ;
        RECT 81.025 134.215 81.195 134.385 ;
        RECT 81.485 134.215 81.655 134.385 ;
        RECT 81.945 134.215 82.115 134.385 ;
        RECT 82.405 134.215 82.575 134.385 ;
        RECT 82.865 134.215 83.035 134.385 ;
        RECT 83.325 134.215 83.495 134.385 ;
        RECT 83.785 134.215 83.955 134.385 ;
        RECT 84.245 134.215 84.415 134.385 ;
        RECT 84.705 134.215 84.875 134.385 ;
        RECT 85.165 134.215 85.335 134.385 ;
        RECT 85.625 134.215 85.795 134.385 ;
        RECT 86.085 134.215 86.255 134.385 ;
        RECT 86.545 134.215 86.715 134.385 ;
        RECT 87.005 134.215 87.175 134.385 ;
        RECT 87.465 134.215 87.635 134.385 ;
        RECT 87.925 134.215 88.095 134.385 ;
        RECT 88.385 134.215 88.555 134.385 ;
        RECT 88.845 134.215 89.015 134.385 ;
        RECT 89.305 134.215 89.475 134.385 ;
        RECT 89.765 134.215 89.935 134.385 ;
        RECT 90.225 134.215 90.395 134.385 ;
        RECT 90.685 134.215 90.855 134.385 ;
        RECT 91.145 134.215 91.315 134.385 ;
        RECT 91.605 134.215 91.775 134.385 ;
        RECT 92.065 134.215 92.235 134.385 ;
        RECT 92.525 134.215 92.695 134.385 ;
        RECT 92.985 134.215 93.155 134.385 ;
        RECT 93.445 134.215 93.615 134.385 ;
        RECT 93.905 134.215 94.075 134.385 ;
        RECT 94.365 134.215 94.535 134.385 ;
        RECT 94.825 134.215 94.995 134.385 ;
        RECT 95.285 134.215 95.455 134.385 ;
        RECT 95.745 134.215 95.915 134.385 ;
        RECT 96.205 134.215 96.375 134.385 ;
        RECT 96.665 134.215 96.835 134.385 ;
        RECT 97.125 134.215 97.295 134.385 ;
        RECT 97.585 134.215 97.755 134.385 ;
        RECT 98.045 134.215 98.215 134.385 ;
        RECT 98.505 134.215 98.675 134.385 ;
        RECT 98.965 134.215 99.135 134.385 ;
        RECT 99.425 134.215 99.595 134.385 ;
        RECT 99.885 134.215 100.055 134.385 ;
        RECT 100.345 134.215 100.515 134.385 ;
        RECT 100.805 134.215 100.975 134.385 ;
        RECT 101.265 134.215 101.435 134.385 ;
        RECT 101.725 134.215 101.895 134.385 ;
        RECT 102.185 134.215 102.355 134.385 ;
        RECT 102.645 134.215 102.815 134.385 ;
        RECT 103.105 134.215 103.275 134.385 ;
        RECT 103.565 134.215 103.735 134.385 ;
        RECT 104.025 134.215 104.195 134.385 ;
        RECT 104.485 134.215 104.655 134.385 ;
        RECT 104.945 134.215 105.115 134.385 ;
        RECT 105.405 134.215 105.575 134.385 ;
        RECT 105.865 134.215 106.035 134.385 ;
        RECT 106.325 134.215 106.495 134.385 ;
        RECT 106.785 134.215 106.955 134.385 ;
        RECT 107.245 134.215 107.415 134.385 ;
        RECT 107.705 134.215 107.875 134.385 ;
        RECT 108.165 134.215 108.335 134.385 ;
        RECT 108.625 134.215 108.795 134.385 ;
        RECT 109.085 134.215 109.255 134.385 ;
        RECT 109.545 134.215 109.715 134.385 ;
        RECT 110.005 134.215 110.175 134.385 ;
        RECT 110.465 134.215 110.635 134.385 ;
        RECT 110.925 134.215 111.095 134.385 ;
        RECT 111.385 134.215 111.555 134.385 ;
        RECT 111.845 134.215 112.015 134.385 ;
        RECT 112.305 134.215 112.475 134.385 ;
        RECT 112.765 134.215 112.935 134.385 ;
        RECT 113.225 134.215 113.395 134.385 ;
        RECT 113.685 134.215 113.855 134.385 ;
        RECT 114.145 134.215 114.315 134.385 ;
        RECT 114.605 134.215 114.775 134.385 ;
        RECT 115.065 134.215 115.235 134.385 ;
        RECT 115.525 134.215 115.695 134.385 ;
        RECT 115.985 134.215 116.155 134.385 ;
        RECT 116.445 134.215 116.615 134.385 ;
        RECT 116.905 134.215 117.075 134.385 ;
        RECT 117.365 134.215 117.535 134.385 ;
        RECT 117.825 134.215 117.995 134.385 ;
        RECT 118.285 134.215 118.455 134.385 ;
        RECT 118.745 134.215 118.915 134.385 ;
        RECT 119.205 134.215 119.375 134.385 ;
        RECT 119.665 134.215 119.835 134.385 ;
        RECT 120.125 134.215 120.295 134.385 ;
        RECT 120.585 134.215 120.755 134.385 ;
        RECT 121.045 134.215 121.215 134.385 ;
        RECT 121.505 134.215 121.675 134.385 ;
        RECT 121.965 134.215 122.135 134.385 ;
        RECT 122.425 134.215 122.595 134.385 ;
        RECT 122.885 134.215 123.055 134.385 ;
        RECT 123.345 134.215 123.515 134.385 ;
        RECT 123.805 134.215 123.975 134.385 ;
        RECT 124.265 134.215 124.435 134.385 ;
        RECT 124.725 134.215 124.895 134.385 ;
        RECT 125.185 134.215 125.355 134.385 ;
        RECT 125.645 134.215 125.815 134.385 ;
        RECT 126.105 134.215 126.275 134.385 ;
        RECT 126.565 134.215 126.735 134.385 ;
        RECT 127.025 134.215 127.195 134.385 ;
        RECT 127.485 134.215 127.655 134.385 ;
        RECT 127.945 134.215 128.115 134.385 ;
        RECT 128.405 134.215 128.575 134.385 ;
        RECT 128.865 134.215 129.035 134.385 ;
        RECT 129.325 134.215 129.495 134.385 ;
        RECT 129.785 134.215 129.955 134.385 ;
        RECT 130.245 134.215 130.415 134.385 ;
        RECT 130.705 134.215 130.875 134.385 ;
        RECT 131.165 134.215 131.335 134.385 ;
        RECT 131.625 134.215 131.795 134.385 ;
        RECT 132.085 134.215 132.255 134.385 ;
        RECT 132.545 134.215 132.715 134.385 ;
        RECT 133.005 134.215 133.175 134.385 ;
        RECT 133.465 134.215 133.635 134.385 ;
        RECT 133.925 134.215 134.095 134.385 ;
        RECT 134.385 134.215 134.555 134.385 ;
        RECT 134.845 134.215 135.015 134.385 ;
        RECT 135.305 134.215 135.475 134.385 ;
        RECT 135.765 134.215 135.935 134.385 ;
        RECT 136.225 134.215 136.395 134.385 ;
        RECT 136.685 134.215 136.855 134.385 ;
        RECT 137.145 134.215 137.315 134.385 ;
        RECT 137.605 134.215 137.775 134.385 ;
        RECT 138.065 134.215 138.235 134.385 ;
        RECT 138.525 134.215 138.695 134.385 ;
        RECT 138.985 134.215 139.155 134.385 ;
        RECT 50.665 131.495 50.835 131.665 ;
        RECT 51.125 131.495 51.295 131.665 ;
        RECT 51.585 131.495 51.755 131.665 ;
        RECT 52.045 131.495 52.215 131.665 ;
        RECT 52.505 131.495 52.675 131.665 ;
        RECT 52.965 131.495 53.135 131.665 ;
        RECT 53.425 131.495 53.595 131.665 ;
        RECT 53.885 131.495 54.055 131.665 ;
        RECT 54.345 131.495 54.515 131.665 ;
        RECT 54.805 131.495 54.975 131.665 ;
        RECT 55.265 131.495 55.435 131.665 ;
        RECT 55.725 131.495 55.895 131.665 ;
        RECT 56.185 131.495 56.355 131.665 ;
        RECT 56.645 131.495 56.815 131.665 ;
        RECT 57.105 131.495 57.275 131.665 ;
        RECT 57.565 131.495 57.735 131.665 ;
        RECT 58.025 131.495 58.195 131.665 ;
        RECT 58.485 131.495 58.655 131.665 ;
        RECT 58.945 131.495 59.115 131.665 ;
        RECT 59.405 131.495 59.575 131.665 ;
        RECT 59.865 131.495 60.035 131.665 ;
        RECT 60.325 131.495 60.495 131.665 ;
        RECT 60.785 131.495 60.955 131.665 ;
        RECT 61.245 131.495 61.415 131.665 ;
        RECT 61.705 131.495 61.875 131.665 ;
        RECT 62.165 131.495 62.335 131.665 ;
        RECT 62.625 131.495 62.795 131.665 ;
        RECT 63.085 131.495 63.255 131.665 ;
        RECT 63.545 131.495 63.715 131.665 ;
        RECT 64.005 131.495 64.175 131.665 ;
        RECT 64.465 131.495 64.635 131.665 ;
        RECT 64.925 131.495 65.095 131.665 ;
        RECT 65.385 131.495 65.555 131.665 ;
        RECT 65.845 131.495 66.015 131.665 ;
        RECT 66.305 131.495 66.475 131.665 ;
        RECT 66.765 131.495 66.935 131.665 ;
        RECT 67.225 131.495 67.395 131.665 ;
        RECT 67.685 131.495 67.855 131.665 ;
        RECT 68.145 131.495 68.315 131.665 ;
        RECT 68.605 131.495 68.775 131.665 ;
        RECT 69.065 131.495 69.235 131.665 ;
        RECT 69.525 131.495 69.695 131.665 ;
        RECT 69.985 131.495 70.155 131.665 ;
        RECT 70.445 131.495 70.615 131.665 ;
        RECT 70.905 131.495 71.075 131.665 ;
        RECT 71.365 131.495 71.535 131.665 ;
        RECT 71.825 131.495 71.995 131.665 ;
        RECT 72.285 131.495 72.455 131.665 ;
        RECT 72.745 131.495 72.915 131.665 ;
        RECT 73.205 131.495 73.375 131.665 ;
        RECT 73.665 131.495 73.835 131.665 ;
        RECT 74.125 131.495 74.295 131.665 ;
        RECT 74.585 131.495 74.755 131.665 ;
        RECT 75.045 131.495 75.215 131.665 ;
        RECT 75.505 131.495 75.675 131.665 ;
        RECT 75.965 131.495 76.135 131.665 ;
        RECT 76.425 131.495 76.595 131.665 ;
        RECT 76.885 131.495 77.055 131.665 ;
        RECT 77.345 131.495 77.515 131.665 ;
        RECT 77.805 131.495 77.975 131.665 ;
        RECT 78.265 131.495 78.435 131.665 ;
        RECT 78.725 131.495 78.895 131.665 ;
        RECT 79.185 131.495 79.355 131.665 ;
        RECT 79.645 131.495 79.815 131.665 ;
        RECT 80.105 131.495 80.275 131.665 ;
        RECT 80.565 131.495 80.735 131.665 ;
        RECT 81.025 131.495 81.195 131.665 ;
        RECT 81.485 131.495 81.655 131.665 ;
        RECT 81.945 131.495 82.115 131.665 ;
        RECT 82.405 131.495 82.575 131.665 ;
        RECT 82.865 131.495 83.035 131.665 ;
        RECT 83.325 131.495 83.495 131.665 ;
        RECT 83.785 131.495 83.955 131.665 ;
        RECT 84.245 131.495 84.415 131.665 ;
        RECT 84.705 131.495 84.875 131.665 ;
        RECT 85.165 131.495 85.335 131.665 ;
        RECT 85.625 131.495 85.795 131.665 ;
        RECT 86.085 131.495 86.255 131.665 ;
        RECT 86.545 131.495 86.715 131.665 ;
        RECT 87.005 131.495 87.175 131.665 ;
        RECT 87.465 131.495 87.635 131.665 ;
        RECT 87.925 131.495 88.095 131.665 ;
        RECT 88.385 131.495 88.555 131.665 ;
        RECT 88.845 131.495 89.015 131.665 ;
        RECT 89.305 131.495 89.475 131.665 ;
        RECT 89.765 131.495 89.935 131.665 ;
        RECT 90.225 131.495 90.395 131.665 ;
        RECT 90.685 131.495 90.855 131.665 ;
        RECT 91.145 131.495 91.315 131.665 ;
        RECT 91.605 131.495 91.775 131.665 ;
        RECT 92.065 131.495 92.235 131.665 ;
        RECT 92.525 131.495 92.695 131.665 ;
        RECT 92.985 131.495 93.155 131.665 ;
        RECT 93.445 131.495 93.615 131.665 ;
        RECT 93.905 131.495 94.075 131.665 ;
        RECT 94.365 131.495 94.535 131.665 ;
        RECT 94.825 131.495 94.995 131.665 ;
        RECT 95.285 131.495 95.455 131.665 ;
        RECT 95.745 131.495 95.915 131.665 ;
        RECT 96.205 131.495 96.375 131.665 ;
        RECT 96.665 131.495 96.835 131.665 ;
        RECT 97.125 131.495 97.295 131.665 ;
        RECT 97.585 131.495 97.755 131.665 ;
        RECT 98.045 131.495 98.215 131.665 ;
        RECT 98.505 131.495 98.675 131.665 ;
        RECT 98.965 131.495 99.135 131.665 ;
        RECT 99.425 131.495 99.595 131.665 ;
        RECT 99.885 131.495 100.055 131.665 ;
        RECT 100.345 131.495 100.515 131.665 ;
        RECT 100.805 131.495 100.975 131.665 ;
        RECT 101.265 131.495 101.435 131.665 ;
        RECT 101.725 131.495 101.895 131.665 ;
        RECT 102.185 131.495 102.355 131.665 ;
        RECT 102.645 131.495 102.815 131.665 ;
        RECT 103.105 131.495 103.275 131.665 ;
        RECT 103.565 131.495 103.735 131.665 ;
        RECT 104.025 131.495 104.195 131.665 ;
        RECT 104.485 131.495 104.655 131.665 ;
        RECT 104.945 131.495 105.115 131.665 ;
        RECT 105.405 131.495 105.575 131.665 ;
        RECT 105.865 131.495 106.035 131.665 ;
        RECT 106.325 131.495 106.495 131.665 ;
        RECT 106.785 131.495 106.955 131.665 ;
        RECT 107.245 131.495 107.415 131.665 ;
        RECT 107.705 131.495 107.875 131.665 ;
        RECT 108.165 131.495 108.335 131.665 ;
        RECT 108.625 131.495 108.795 131.665 ;
        RECT 109.085 131.495 109.255 131.665 ;
        RECT 109.545 131.495 109.715 131.665 ;
        RECT 110.005 131.495 110.175 131.665 ;
        RECT 110.465 131.495 110.635 131.665 ;
        RECT 110.925 131.495 111.095 131.665 ;
        RECT 111.385 131.495 111.555 131.665 ;
        RECT 111.845 131.495 112.015 131.665 ;
        RECT 112.305 131.495 112.475 131.665 ;
        RECT 112.765 131.495 112.935 131.665 ;
        RECT 113.225 131.495 113.395 131.665 ;
        RECT 113.685 131.495 113.855 131.665 ;
        RECT 114.145 131.495 114.315 131.665 ;
        RECT 114.605 131.495 114.775 131.665 ;
        RECT 115.065 131.495 115.235 131.665 ;
        RECT 115.525 131.495 115.695 131.665 ;
        RECT 115.985 131.495 116.155 131.665 ;
        RECT 116.445 131.495 116.615 131.665 ;
        RECT 116.905 131.495 117.075 131.665 ;
        RECT 117.365 131.495 117.535 131.665 ;
        RECT 117.825 131.495 117.995 131.665 ;
        RECT 118.285 131.495 118.455 131.665 ;
        RECT 118.745 131.495 118.915 131.665 ;
        RECT 119.205 131.495 119.375 131.665 ;
        RECT 119.665 131.495 119.835 131.665 ;
        RECT 120.125 131.495 120.295 131.665 ;
        RECT 120.585 131.495 120.755 131.665 ;
        RECT 121.045 131.495 121.215 131.665 ;
        RECT 121.505 131.495 121.675 131.665 ;
        RECT 121.965 131.495 122.135 131.665 ;
        RECT 122.425 131.495 122.595 131.665 ;
        RECT 122.885 131.495 123.055 131.665 ;
        RECT 123.345 131.495 123.515 131.665 ;
        RECT 123.805 131.495 123.975 131.665 ;
        RECT 124.265 131.495 124.435 131.665 ;
        RECT 124.725 131.495 124.895 131.665 ;
        RECT 125.185 131.495 125.355 131.665 ;
        RECT 125.645 131.495 125.815 131.665 ;
        RECT 126.105 131.495 126.275 131.665 ;
        RECT 126.565 131.495 126.735 131.665 ;
        RECT 127.025 131.495 127.195 131.665 ;
        RECT 127.485 131.495 127.655 131.665 ;
        RECT 127.945 131.495 128.115 131.665 ;
        RECT 128.405 131.495 128.575 131.665 ;
        RECT 128.865 131.495 129.035 131.665 ;
        RECT 129.325 131.495 129.495 131.665 ;
        RECT 129.785 131.495 129.955 131.665 ;
        RECT 130.245 131.495 130.415 131.665 ;
        RECT 130.705 131.495 130.875 131.665 ;
        RECT 131.165 131.495 131.335 131.665 ;
        RECT 131.625 131.495 131.795 131.665 ;
        RECT 132.085 131.495 132.255 131.665 ;
        RECT 132.545 131.495 132.715 131.665 ;
        RECT 133.005 131.495 133.175 131.665 ;
        RECT 133.465 131.495 133.635 131.665 ;
        RECT 133.925 131.495 134.095 131.665 ;
        RECT 134.385 131.495 134.555 131.665 ;
        RECT 134.845 131.495 135.015 131.665 ;
        RECT 135.305 131.495 135.475 131.665 ;
        RECT 135.765 131.495 135.935 131.665 ;
        RECT 136.225 131.495 136.395 131.665 ;
        RECT 136.685 131.495 136.855 131.665 ;
        RECT 137.145 131.495 137.315 131.665 ;
        RECT 137.605 131.495 137.775 131.665 ;
        RECT 138.065 131.495 138.235 131.665 ;
        RECT 138.525 131.495 138.695 131.665 ;
        RECT 138.985 131.495 139.155 131.665 ;
        RECT 50.665 128.775 50.835 128.945 ;
        RECT 51.125 128.775 51.295 128.945 ;
        RECT 51.585 128.775 51.755 128.945 ;
        RECT 52.045 128.775 52.215 128.945 ;
        RECT 52.505 128.775 52.675 128.945 ;
        RECT 52.965 128.775 53.135 128.945 ;
        RECT 53.425 128.775 53.595 128.945 ;
        RECT 53.885 128.775 54.055 128.945 ;
        RECT 54.345 128.775 54.515 128.945 ;
        RECT 54.805 128.775 54.975 128.945 ;
        RECT 55.265 128.775 55.435 128.945 ;
        RECT 55.725 128.775 55.895 128.945 ;
        RECT 56.185 128.775 56.355 128.945 ;
        RECT 56.645 128.775 56.815 128.945 ;
        RECT 57.105 128.775 57.275 128.945 ;
        RECT 57.565 128.775 57.735 128.945 ;
        RECT 58.025 128.775 58.195 128.945 ;
        RECT 58.485 128.775 58.655 128.945 ;
        RECT 58.945 128.775 59.115 128.945 ;
        RECT 59.405 128.775 59.575 128.945 ;
        RECT 59.865 128.775 60.035 128.945 ;
        RECT 60.325 128.775 60.495 128.945 ;
        RECT 60.785 128.775 60.955 128.945 ;
        RECT 61.245 128.775 61.415 128.945 ;
        RECT 61.705 128.775 61.875 128.945 ;
        RECT 62.165 128.775 62.335 128.945 ;
        RECT 62.625 128.775 62.795 128.945 ;
        RECT 63.085 128.775 63.255 128.945 ;
        RECT 63.545 128.775 63.715 128.945 ;
        RECT 64.005 128.775 64.175 128.945 ;
        RECT 64.465 128.775 64.635 128.945 ;
        RECT 64.925 128.775 65.095 128.945 ;
        RECT 65.385 128.775 65.555 128.945 ;
        RECT 65.845 128.775 66.015 128.945 ;
        RECT 66.305 128.775 66.475 128.945 ;
        RECT 66.765 128.775 66.935 128.945 ;
        RECT 67.225 128.775 67.395 128.945 ;
        RECT 67.685 128.775 67.855 128.945 ;
        RECT 68.145 128.775 68.315 128.945 ;
        RECT 68.605 128.775 68.775 128.945 ;
        RECT 69.065 128.775 69.235 128.945 ;
        RECT 69.525 128.775 69.695 128.945 ;
        RECT 69.985 128.775 70.155 128.945 ;
        RECT 70.445 128.775 70.615 128.945 ;
        RECT 70.905 128.775 71.075 128.945 ;
        RECT 71.365 128.775 71.535 128.945 ;
        RECT 71.825 128.775 71.995 128.945 ;
        RECT 72.285 128.775 72.455 128.945 ;
        RECT 72.745 128.775 72.915 128.945 ;
        RECT 73.205 128.775 73.375 128.945 ;
        RECT 73.665 128.775 73.835 128.945 ;
        RECT 74.125 128.775 74.295 128.945 ;
        RECT 74.585 128.775 74.755 128.945 ;
        RECT 75.045 128.775 75.215 128.945 ;
        RECT 75.505 128.775 75.675 128.945 ;
        RECT 75.965 128.775 76.135 128.945 ;
        RECT 76.425 128.775 76.595 128.945 ;
        RECT 76.885 128.775 77.055 128.945 ;
        RECT 77.345 128.775 77.515 128.945 ;
        RECT 77.805 128.775 77.975 128.945 ;
        RECT 78.265 128.775 78.435 128.945 ;
        RECT 78.725 128.775 78.895 128.945 ;
        RECT 79.185 128.775 79.355 128.945 ;
        RECT 79.645 128.775 79.815 128.945 ;
        RECT 80.105 128.775 80.275 128.945 ;
        RECT 80.565 128.775 80.735 128.945 ;
        RECT 81.025 128.775 81.195 128.945 ;
        RECT 81.485 128.775 81.655 128.945 ;
        RECT 81.945 128.775 82.115 128.945 ;
        RECT 82.405 128.775 82.575 128.945 ;
        RECT 82.865 128.775 83.035 128.945 ;
        RECT 83.325 128.775 83.495 128.945 ;
        RECT 83.785 128.775 83.955 128.945 ;
        RECT 84.245 128.775 84.415 128.945 ;
        RECT 84.705 128.775 84.875 128.945 ;
        RECT 85.165 128.775 85.335 128.945 ;
        RECT 85.625 128.775 85.795 128.945 ;
        RECT 86.085 128.775 86.255 128.945 ;
        RECT 86.545 128.775 86.715 128.945 ;
        RECT 87.005 128.775 87.175 128.945 ;
        RECT 87.465 128.775 87.635 128.945 ;
        RECT 87.925 128.775 88.095 128.945 ;
        RECT 88.385 128.775 88.555 128.945 ;
        RECT 88.845 128.775 89.015 128.945 ;
        RECT 89.305 128.775 89.475 128.945 ;
        RECT 89.765 128.775 89.935 128.945 ;
        RECT 90.225 128.775 90.395 128.945 ;
        RECT 90.685 128.775 90.855 128.945 ;
        RECT 91.145 128.775 91.315 128.945 ;
        RECT 91.605 128.775 91.775 128.945 ;
        RECT 92.065 128.775 92.235 128.945 ;
        RECT 92.525 128.775 92.695 128.945 ;
        RECT 92.985 128.775 93.155 128.945 ;
        RECT 93.445 128.775 93.615 128.945 ;
        RECT 93.905 128.775 94.075 128.945 ;
        RECT 94.365 128.775 94.535 128.945 ;
        RECT 94.825 128.775 94.995 128.945 ;
        RECT 95.285 128.775 95.455 128.945 ;
        RECT 95.745 128.775 95.915 128.945 ;
        RECT 96.205 128.775 96.375 128.945 ;
        RECT 96.665 128.775 96.835 128.945 ;
        RECT 97.125 128.775 97.295 128.945 ;
        RECT 97.585 128.775 97.755 128.945 ;
        RECT 98.045 128.775 98.215 128.945 ;
        RECT 98.505 128.775 98.675 128.945 ;
        RECT 98.965 128.775 99.135 128.945 ;
        RECT 99.425 128.775 99.595 128.945 ;
        RECT 99.885 128.775 100.055 128.945 ;
        RECT 100.345 128.775 100.515 128.945 ;
        RECT 100.805 128.775 100.975 128.945 ;
        RECT 101.265 128.775 101.435 128.945 ;
        RECT 101.725 128.775 101.895 128.945 ;
        RECT 102.185 128.775 102.355 128.945 ;
        RECT 102.645 128.775 102.815 128.945 ;
        RECT 103.105 128.775 103.275 128.945 ;
        RECT 103.565 128.775 103.735 128.945 ;
        RECT 104.025 128.775 104.195 128.945 ;
        RECT 104.485 128.775 104.655 128.945 ;
        RECT 104.945 128.775 105.115 128.945 ;
        RECT 105.405 128.775 105.575 128.945 ;
        RECT 105.865 128.775 106.035 128.945 ;
        RECT 106.325 128.775 106.495 128.945 ;
        RECT 106.785 128.775 106.955 128.945 ;
        RECT 107.245 128.775 107.415 128.945 ;
        RECT 107.705 128.775 107.875 128.945 ;
        RECT 108.165 128.775 108.335 128.945 ;
        RECT 108.625 128.775 108.795 128.945 ;
        RECT 109.085 128.775 109.255 128.945 ;
        RECT 109.545 128.775 109.715 128.945 ;
        RECT 110.005 128.775 110.175 128.945 ;
        RECT 110.465 128.775 110.635 128.945 ;
        RECT 110.925 128.775 111.095 128.945 ;
        RECT 111.385 128.775 111.555 128.945 ;
        RECT 111.845 128.775 112.015 128.945 ;
        RECT 112.305 128.775 112.475 128.945 ;
        RECT 112.765 128.775 112.935 128.945 ;
        RECT 113.225 128.775 113.395 128.945 ;
        RECT 113.685 128.775 113.855 128.945 ;
        RECT 114.145 128.775 114.315 128.945 ;
        RECT 114.605 128.775 114.775 128.945 ;
        RECT 115.065 128.775 115.235 128.945 ;
        RECT 115.525 128.775 115.695 128.945 ;
        RECT 115.985 128.775 116.155 128.945 ;
        RECT 116.445 128.775 116.615 128.945 ;
        RECT 116.905 128.775 117.075 128.945 ;
        RECT 117.365 128.775 117.535 128.945 ;
        RECT 117.825 128.775 117.995 128.945 ;
        RECT 118.285 128.775 118.455 128.945 ;
        RECT 118.745 128.775 118.915 128.945 ;
        RECT 119.205 128.775 119.375 128.945 ;
        RECT 119.665 128.775 119.835 128.945 ;
        RECT 120.125 128.775 120.295 128.945 ;
        RECT 120.585 128.775 120.755 128.945 ;
        RECT 121.045 128.775 121.215 128.945 ;
        RECT 121.505 128.775 121.675 128.945 ;
        RECT 121.965 128.775 122.135 128.945 ;
        RECT 122.425 128.775 122.595 128.945 ;
        RECT 122.885 128.775 123.055 128.945 ;
        RECT 123.345 128.775 123.515 128.945 ;
        RECT 123.805 128.775 123.975 128.945 ;
        RECT 124.265 128.775 124.435 128.945 ;
        RECT 124.725 128.775 124.895 128.945 ;
        RECT 125.185 128.775 125.355 128.945 ;
        RECT 125.645 128.775 125.815 128.945 ;
        RECT 126.105 128.775 126.275 128.945 ;
        RECT 126.565 128.775 126.735 128.945 ;
        RECT 127.025 128.775 127.195 128.945 ;
        RECT 127.485 128.775 127.655 128.945 ;
        RECT 127.945 128.775 128.115 128.945 ;
        RECT 128.405 128.775 128.575 128.945 ;
        RECT 128.865 128.775 129.035 128.945 ;
        RECT 129.325 128.775 129.495 128.945 ;
        RECT 129.785 128.775 129.955 128.945 ;
        RECT 130.245 128.775 130.415 128.945 ;
        RECT 130.705 128.775 130.875 128.945 ;
        RECT 131.165 128.775 131.335 128.945 ;
        RECT 131.625 128.775 131.795 128.945 ;
        RECT 132.085 128.775 132.255 128.945 ;
        RECT 132.545 128.775 132.715 128.945 ;
        RECT 133.005 128.775 133.175 128.945 ;
        RECT 133.465 128.775 133.635 128.945 ;
        RECT 133.925 128.775 134.095 128.945 ;
        RECT 134.385 128.775 134.555 128.945 ;
        RECT 134.845 128.775 135.015 128.945 ;
        RECT 135.305 128.775 135.475 128.945 ;
        RECT 135.765 128.775 135.935 128.945 ;
        RECT 136.225 128.775 136.395 128.945 ;
        RECT 136.685 128.775 136.855 128.945 ;
        RECT 137.145 128.775 137.315 128.945 ;
        RECT 137.605 128.775 137.775 128.945 ;
        RECT 138.065 128.775 138.235 128.945 ;
        RECT 138.525 128.775 138.695 128.945 ;
        RECT 138.985 128.775 139.155 128.945 ;
        RECT 50.665 126.055 50.835 126.225 ;
        RECT 51.125 126.055 51.295 126.225 ;
        RECT 51.585 126.055 51.755 126.225 ;
        RECT 52.045 126.055 52.215 126.225 ;
        RECT 52.505 126.055 52.675 126.225 ;
        RECT 52.965 126.055 53.135 126.225 ;
        RECT 53.425 126.055 53.595 126.225 ;
        RECT 53.885 126.055 54.055 126.225 ;
        RECT 54.345 126.055 54.515 126.225 ;
        RECT 54.805 126.055 54.975 126.225 ;
        RECT 55.265 126.055 55.435 126.225 ;
        RECT 55.725 126.055 55.895 126.225 ;
        RECT 56.185 126.055 56.355 126.225 ;
        RECT 56.645 126.055 56.815 126.225 ;
        RECT 57.105 126.055 57.275 126.225 ;
        RECT 57.565 126.055 57.735 126.225 ;
        RECT 58.025 126.055 58.195 126.225 ;
        RECT 58.485 126.055 58.655 126.225 ;
        RECT 58.945 126.055 59.115 126.225 ;
        RECT 59.405 126.055 59.575 126.225 ;
        RECT 59.865 126.055 60.035 126.225 ;
        RECT 60.325 126.055 60.495 126.225 ;
        RECT 60.785 126.055 60.955 126.225 ;
        RECT 61.245 126.055 61.415 126.225 ;
        RECT 61.705 126.055 61.875 126.225 ;
        RECT 62.165 126.055 62.335 126.225 ;
        RECT 62.625 126.055 62.795 126.225 ;
        RECT 63.085 126.055 63.255 126.225 ;
        RECT 63.545 126.055 63.715 126.225 ;
        RECT 64.005 126.055 64.175 126.225 ;
        RECT 64.465 126.055 64.635 126.225 ;
        RECT 64.925 126.055 65.095 126.225 ;
        RECT 65.385 126.055 65.555 126.225 ;
        RECT 65.845 126.055 66.015 126.225 ;
        RECT 66.305 126.055 66.475 126.225 ;
        RECT 66.765 126.055 66.935 126.225 ;
        RECT 67.225 126.055 67.395 126.225 ;
        RECT 67.685 126.055 67.855 126.225 ;
        RECT 68.145 126.055 68.315 126.225 ;
        RECT 68.605 126.055 68.775 126.225 ;
        RECT 69.065 126.055 69.235 126.225 ;
        RECT 69.525 126.055 69.695 126.225 ;
        RECT 69.985 126.055 70.155 126.225 ;
        RECT 70.445 126.055 70.615 126.225 ;
        RECT 70.905 126.055 71.075 126.225 ;
        RECT 71.365 126.055 71.535 126.225 ;
        RECT 71.825 126.055 71.995 126.225 ;
        RECT 72.285 126.055 72.455 126.225 ;
        RECT 72.745 126.055 72.915 126.225 ;
        RECT 73.205 126.055 73.375 126.225 ;
        RECT 73.665 126.055 73.835 126.225 ;
        RECT 74.125 126.055 74.295 126.225 ;
        RECT 74.585 126.055 74.755 126.225 ;
        RECT 75.045 126.055 75.215 126.225 ;
        RECT 75.505 126.055 75.675 126.225 ;
        RECT 75.965 126.055 76.135 126.225 ;
        RECT 76.425 126.055 76.595 126.225 ;
        RECT 76.885 126.055 77.055 126.225 ;
        RECT 77.345 126.055 77.515 126.225 ;
        RECT 77.805 126.055 77.975 126.225 ;
        RECT 78.265 126.055 78.435 126.225 ;
        RECT 78.725 126.055 78.895 126.225 ;
        RECT 79.185 126.055 79.355 126.225 ;
        RECT 79.645 126.055 79.815 126.225 ;
        RECT 80.105 126.055 80.275 126.225 ;
        RECT 80.565 126.055 80.735 126.225 ;
        RECT 81.025 126.055 81.195 126.225 ;
        RECT 81.485 126.055 81.655 126.225 ;
        RECT 81.945 126.055 82.115 126.225 ;
        RECT 82.405 126.055 82.575 126.225 ;
        RECT 82.865 126.055 83.035 126.225 ;
        RECT 83.325 126.055 83.495 126.225 ;
        RECT 83.785 126.055 83.955 126.225 ;
        RECT 84.245 126.055 84.415 126.225 ;
        RECT 84.705 126.055 84.875 126.225 ;
        RECT 85.165 126.055 85.335 126.225 ;
        RECT 85.625 126.055 85.795 126.225 ;
        RECT 86.085 126.055 86.255 126.225 ;
        RECT 86.545 126.055 86.715 126.225 ;
        RECT 87.005 126.055 87.175 126.225 ;
        RECT 87.465 126.055 87.635 126.225 ;
        RECT 87.925 126.055 88.095 126.225 ;
        RECT 88.385 126.055 88.555 126.225 ;
        RECT 88.845 126.055 89.015 126.225 ;
        RECT 89.305 126.055 89.475 126.225 ;
        RECT 89.765 126.055 89.935 126.225 ;
        RECT 90.225 126.055 90.395 126.225 ;
        RECT 90.685 126.055 90.855 126.225 ;
        RECT 91.145 126.055 91.315 126.225 ;
        RECT 91.605 126.055 91.775 126.225 ;
        RECT 92.065 126.055 92.235 126.225 ;
        RECT 92.525 126.055 92.695 126.225 ;
        RECT 92.985 126.055 93.155 126.225 ;
        RECT 93.445 126.055 93.615 126.225 ;
        RECT 93.905 126.055 94.075 126.225 ;
        RECT 94.365 126.055 94.535 126.225 ;
        RECT 94.825 126.055 94.995 126.225 ;
        RECT 95.285 126.055 95.455 126.225 ;
        RECT 95.745 126.055 95.915 126.225 ;
        RECT 96.205 126.055 96.375 126.225 ;
        RECT 96.665 126.055 96.835 126.225 ;
        RECT 97.125 126.055 97.295 126.225 ;
        RECT 97.585 126.055 97.755 126.225 ;
        RECT 98.045 126.055 98.215 126.225 ;
        RECT 98.505 126.055 98.675 126.225 ;
        RECT 98.965 126.055 99.135 126.225 ;
        RECT 99.425 126.055 99.595 126.225 ;
        RECT 99.885 126.055 100.055 126.225 ;
        RECT 100.345 126.055 100.515 126.225 ;
        RECT 100.805 126.055 100.975 126.225 ;
        RECT 101.265 126.055 101.435 126.225 ;
        RECT 101.725 126.055 101.895 126.225 ;
        RECT 102.185 126.055 102.355 126.225 ;
        RECT 102.645 126.055 102.815 126.225 ;
        RECT 103.105 126.055 103.275 126.225 ;
        RECT 103.565 126.055 103.735 126.225 ;
        RECT 104.025 126.055 104.195 126.225 ;
        RECT 104.485 126.055 104.655 126.225 ;
        RECT 104.945 126.055 105.115 126.225 ;
        RECT 105.405 126.055 105.575 126.225 ;
        RECT 105.865 126.055 106.035 126.225 ;
        RECT 106.325 126.055 106.495 126.225 ;
        RECT 106.785 126.055 106.955 126.225 ;
        RECT 107.245 126.055 107.415 126.225 ;
        RECT 107.705 126.055 107.875 126.225 ;
        RECT 108.165 126.055 108.335 126.225 ;
        RECT 108.625 126.055 108.795 126.225 ;
        RECT 109.085 126.055 109.255 126.225 ;
        RECT 109.545 126.055 109.715 126.225 ;
        RECT 110.005 126.055 110.175 126.225 ;
        RECT 110.465 126.055 110.635 126.225 ;
        RECT 110.925 126.055 111.095 126.225 ;
        RECT 111.385 126.055 111.555 126.225 ;
        RECT 111.845 126.055 112.015 126.225 ;
        RECT 112.305 126.055 112.475 126.225 ;
        RECT 112.765 126.055 112.935 126.225 ;
        RECT 113.225 126.055 113.395 126.225 ;
        RECT 113.685 126.055 113.855 126.225 ;
        RECT 114.145 126.055 114.315 126.225 ;
        RECT 114.605 126.055 114.775 126.225 ;
        RECT 115.065 126.055 115.235 126.225 ;
        RECT 115.525 126.055 115.695 126.225 ;
        RECT 115.985 126.055 116.155 126.225 ;
        RECT 116.445 126.055 116.615 126.225 ;
        RECT 116.905 126.055 117.075 126.225 ;
        RECT 117.365 126.055 117.535 126.225 ;
        RECT 117.825 126.055 117.995 126.225 ;
        RECT 118.285 126.055 118.455 126.225 ;
        RECT 118.745 126.055 118.915 126.225 ;
        RECT 119.205 126.055 119.375 126.225 ;
        RECT 119.665 126.055 119.835 126.225 ;
        RECT 120.125 126.055 120.295 126.225 ;
        RECT 120.585 126.055 120.755 126.225 ;
        RECT 121.045 126.055 121.215 126.225 ;
        RECT 121.505 126.055 121.675 126.225 ;
        RECT 121.965 126.055 122.135 126.225 ;
        RECT 122.425 126.055 122.595 126.225 ;
        RECT 122.885 126.055 123.055 126.225 ;
        RECT 123.345 126.055 123.515 126.225 ;
        RECT 123.805 126.055 123.975 126.225 ;
        RECT 124.265 126.055 124.435 126.225 ;
        RECT 124.725 126.055 124.895 126.225 ;
        RECT 125.185 126.055 125.355 126.225 ;
        RECT 125.645 126.055 125.815 126.225 ;
        RECT 126.105 126.055 126.275 126.225 ;
        RECT 126.565 126.055 126.735 126.225 ;
        RECT 127.025 126.055 127.195 126.225 ;
        RECT 127.485 126.055 127.655 126.225 ;
        RECT 127.945 126.055 128.115 126.225 ;
        RECT 128.405 126.055 128.575 126.225 ;
        RECT 128.865 126.055 129.035 126.225 ;
        RECT 129.325 126.055 129.495 126.225 ;
        RECT 129.785 126.055 129.955 126.225 ;
        RECT 130.245 126.055 130.415 126.225 ;
        RECT 130.705 126.055 130.875 126.225 ;
        RECT 131.165 126.055 131.335 126.225 ;
        RECT 131.625 126.055 131.795 126.225 ;
        RECT 132.085 126.055 132.255 126.225 ;
        RECT 132.545 126.055 132.715 126.225 ;
        RECT 133.005 126.055 133.175 126.225 ;
        RECT 133.465 126.055 133.635 126.225 ;
        RECT 133.925 126.055 134.095 126.225 ;
        RECT 134.385 126.055 134.555 126.225 ;
        RECT 134.845 126.055 135.015 126.225 ;
        RECT 135.305 126.055 135.475 126.225 ;
        RECT 135.765 126.055 135.935 126.225 ;
        RECT 136.225 126.055 136.395 126.225 ;
        RECT 136.685 126.055 136.855 126.225 ;
        RECT 137.145 126.055 137.315 126.225 ;
        RECT 137.605 126.055 137.775 126.225 ;
        RECT 138.065 126.055 138.235 126.225 ;
        RECT 138.525 126.055 138.695 126.225 ;
        RECT 138.985 126.055 139.155 126.225 ;
        RECT 50.665 123.335 50.835 123.505 ;
        RECT 51.125 123.335 51.295 123.505 ;
        RECT 51.585 123.335 51.755 123.505 ;
        RECT 52.045 123.335 52.215 123.505 ;
        RECT 52.505 123.335 52.675 123.505 ;
        RECT 52.965 123.335 53.135 123.505 ;
        RECT 53.425 123.335 53.595 123.505 ;
        RECT 53.885 123.335 54.055 123.505 ;
        RECT 54.345 123.335 54.515 123.505 ;
        RECT 54.805 123.335 54.975 123.505 ;
        RECT 55.265 123.335 55.435 123.505 ;
        RECT 55.725 123.335 55.895 123.505 ;
        RECT 56.185 123.335 56.355 123.505 ;
        RECT 56.645 123.335 56.815 123.505 ;
        RECT 57.105 123.335 57.275 123.505 ;
        RECT 57.565 123.335 57.735 123.505 ;
        RECT 58.025 123.335 58.195 123.505 ;
        RECT 58.485 123.335 58.655 123.505 ;
        RECT 58.945 123.335 59.115 123.505 ;
        RECT 59.405 123.335 59.575 123.505 ;
        RECT 59.865 123.335 60.035 123.505 ;
        RECT 60.325 123.335 60.495 123.505 ;
        RECT 60.785 123.335 60.955 123.505 ;
        RECT 61.245 123.335 61.415 123.505 ;
        RECT 61.705 123.335 61.875 123.505 ;
        RECT 62.165 123.335 62.335 123.505 ;
        RECT 62.625 123.335 62.795 123.505 ;
        RECT 63.085 123.335 63.255 123.505 ;
        RECT 63.545 123.335 63.715 123.505 ;
        RECT 64.005 123.335 64.175 123.505 ;
        RECT 64.465 123.335 64.635 123.505 ;
        RECT 64.925 123.335 65.095 123.505 ;
        RECT 65.385 123.335 65.555 123.505 ;
        RECT 65.845 123.335 66.015 123.505 ;
        RECT 66.305 123.335 66.475 123.505 ;
        RECT 66.765 123.335 66.935 123.505 ;
        RECT 67.225 123.335 67.395 123.505 ;
        RECT 67.685 123.335 67.855 123.505 ;
        RECT 68.145 123.335 68.315 123.505 ;
        RECT 68.605 123.335 68.775 123.505 ;
        RECT 69.065 123.335 69.235 123.505 ;
        RECT 69.525 123.335 69.695 123.505 ;
        RECT 69.985 123.335 70.155 123.505 ;
        RECT 70.445 123.335 70.615 123.505 ;
        RECT 70.905 123.335 71.075 123.505 ;
        RECT 71.365 123.335 71.535 123.505 ;
        RECT 71.825 123.335 71.995 123.505 ;
        RECT 72.285 123.335 72.455 123.505 ;
        RECT 72.745 123.335 72.915 123.505 ;
        RECT 73.205 123.335 73.375 123.505 ;
        RECT 73.665 123.335 73.835 123.505 ;
        RECT 74.125 123.335 74.295 123.505 ;
        RECT 74.585 123.335 74.755 123.505 ;
        RECT 75.045 123.335 75.215 123.505 ;
        RECT 75.505 123.335 75.675 123.505 ;
        RECT 75.965 123.335 76.135 123.505 ;
        RECT 76.425 123.335 76.595 123.505 ;
        RECT 76.885 123.335 77.055 123.505 ;
        RECT 77.345 123.335 77.515 123.505 ;
        RECT 77.805 123.335 77.975 123.505 ;
        RECT 78.265 123.335 78.435 123.505 ;
        RECT 78.725 123.335 78.895 123.505 ;
        RECT 79.185 123.335 79.355 123.505 ;
        RECT 79.645 123.335 79.815 123.505 ;
        RECT 80.105 123.335 80.275 123.505 ;
        RECT 80.565 123.335 80.735 123.505 ;
        RECT 81.025 123.335 81.195 123.505 ;
        RECT 81.485 123.335 81.655 123.505 ;
        RECT 81.945 123.335 82.115 123.505 ;
        RECT 82.405 123.335 82.575 123.505 ;
        RECT 82.865 123.335 83.035 123.505 ;
        RECT 83.325 123.335 83.495 123.505 ;
        RECT 83.785 123.335 83.955 123.505 ;
        RECT 84.245 123.335 84.415 123.505 ;
        RECT 84.705 123.335 84.875 123.505 ;
        RECT 85.165 123.335 85.335 123.505 ;
        RECT 85.625 123.335 85.795 123.505 ;
        RECT 86.085 123.335 86.255 123.505 ;
        RECT 86.545 123.335 86.715 123.505 ;
        RECT 87.005 123.335 87.175 123.505 ;
        RECT 87.465 123.335 87.635 123.505 ;
        RECT 87.925 123.335 88.095 123.505 ;
        RECT 88.385 123.335 88.555 123.505 ;
        RECT 88.845 123.335 89.015 123.505 ;
        RECT 89.305 123.335 89.475 123.505 ;
        RECT 89.765 123.335 89.935 123.505 ;
        RECT 90.225 123.335 90.395 123.505 ;
        RECT 90.685 123.335 90.855 123.505 ;
        RECT 91.145 123.335 91.315 123.505 ;
        RECT 91.605 123.335 91.775 123.505 ;
        RECT 92.065 123.335 92.235 123.505 ;
        RECT 92.525 123.335 92.695 123.505 ;
        RECT 92.985 123.335 93.155 123.505 ;
        RECT 93.445 123.335 93.615 123.505 ;
        RECT 93.905 123.335 94.075 123.505 ;
        RECT 94.365 123.335 94.535 123.505 ;
        RECT 94.825 123.335 94.995 123.505 ;
        RECT 95.285 123.335 95.455 123.505 ;
        RECT 95.745 123.335 95.915 123.505 ;
        RECT 96.205 123.335 96.375 123.505 ;
        RECT 96.665 123.335 96.835 123.505 ;
        RECT 97.125 123.335 97.295 123.505 ;
        RECT 97.585 123.335 97.755 123.505 ;
        RECT 98.045 123.335 98.215 123.505 ;
        RECT 98.505 123.335 98.675 123.505 ;
        RECT 98.965 123.335 99.135 123.505 ;
        RECT 99.425 123.335 99.595 123.505 ;
        RECT 99.885 123.335 100.055 123.505 ;
        RECT 100.345 123.335 100.515 123.505 ;
        RECT 100.805 123.335 100.975 123.505 ;
        RECT 101.265 123.335 101.435 123.505 ;
        RECT 101.725 123.335 101.895 123.505 ;
        RECT 102.185 123.335 102.355 123.505 ;
        RECT 102.645 123.335 102.815 123.505 ;
        RECT 103.105 123.335 103.275 123.505 ;
        RECT 103.565 123.335 103.735 123.505 ;
        RECT 104.025 123.335 104.195 123.505 ;
        RECT 104.485 123.335 104.655 123.505 ;
        RECT 104.945 123.335 105.115 123.505 ;
        RECT 105.405 123.335 105.575 123.505 ;
        RECT 105.865 123.335 106.035 123.505 ;
        RECT 106.325 123.335 106.495 123.505 ;
        RECT 106.785 123.335 106.955 123.505 ;
        RECT 107.245 123.335 107.415 123.505 ;
        RECT 107.705 123.335 107.875 123.505 ;
        RECT 108.165 123.335 108.335 123.505 ;
        RECT 108.625 123.335 108.795 123.505 ;
        RECT 109.085 123.335 109.255 123.505 ;
        RECT 109.545 123.335 109.715 123.505 ;
        RECT 110.005 123.335 110.175 123.505 ;
        RECT 110.465 123.335 110.635 123.505 ;
        RECT 110.925 123.335 111.095 123.505 ;
        RECT 111.385 123.335 111.555 123.505 ;
        RECT 111.845 123.335 112.015 123.505 ;
        RECT 112.305 123.335 112.475 123.505 ;
        RECT 112.765 123.335 112.935 123.505 ;
        RECT 113.225 123.335 113.395 123.505 ;
        RECT 113.685 123.335 113.855 123.505 ;
        RECT 114.145 123.335 114.315 123.505 ;
        RECT 114.605 123.335 114.775 123.505 ;
        RECT 115.065 123.335 115.235 123.505 ;
        RECT 115.525 123.335 115.695 123.505 ;
        RECT 115.985 123.335 116.155 123.505 ;
        RECT 116.445 123.335 116.615 123.505 ;
        RECT 116.905 123.335 117.075 123.505 ;
        RECT 117.365 123.335 117.535 123.505 ;
        RECT 117.825 123.335 117.995 123.505 ;
        RECT 118.285 123.335 118.455 123.505 ;
        RECT 118.745 123.335 118.915 123.505 ;
        RECT 119.205 123.335 119.375 123.505 ;
        RECT 119.665 123.335 119.835 123.505 ;
        RECT 120.125 123.335 120.295 123.505 ;
        RECT 120.585 123.335 120.755 123.505 ;
        RECT 121.045 123.335 121.215 123.505 ;
        RECT 121.505 123.335 121.675 123.505 ;
        RECT 121.965 123.335 122.135 123.505 ;
        RECT 122.425 123.335 122.595 123.505 ;
        RECT 122.885 123.335 123.055 123.505 ;
        RECT 123.345 123.335 123.515 123.505 ;
        RECT 123.805 123.335 123.975 123.505 ;
        RECT 124.265 123.335 124.435 123.505 ;
        RECT 124.725 123.335 124.895 123.505 ;
        RECT 125.185 123.335 125.355 123.505 ;
        RECT 125.645 123.335 125.815 123.505 ;
        RECT 126.105 123.335 126.275 123.505 ;
        RECT 126.565 123.335 126.735 123.505 ;
        RECT 127.025 123.335 127.195 123.505 ;
        RECT 127.485 123.335 127.655 123.505 ;
        RECT 127.945 123.335 128.115 123.505 ;
        RECT 128.405 123.335 128.575 123.505 ;
        RECT 128.865 123.335 129.035 123.505 ;
        RECT 129.325 123.335 129.495 123.505 ;
        RECT 129.785 123.335 129.955 123.505 ;
        RECT 130.245 123.335 130.415 123.505 ;
        RECT 130.705 123.335 130.875 123.505 ;
        RECT 131.165 123.335 131.335 123.505 ;
        RECT 131.625 123.335 131.795 123.505 ;
        RECT 132.085 123.335 132.255 123.505 ;
        RECT 132.545 123.335 132.715 123.505 ;
        RECT 133.005 123.335 133.175 123.505 ;
        RECT 133.465 123.335 133.635 123.505 ;
        RECT 133.925 123.335 134.095 123.505 ;
        RECT 134.385 123.335 134.555 123.505 ;
        RECT 134.845 123.335 135.015 123.505 ;
        RECT 135.305 123.335 135.475 123.505 ;
        RECT 135.765 123.335 135.935 123.505 ;
        RECT 136.225 123.335 136.395 123.505 ;
        RECT 136.685 123.335 136.855 123.505 ;
        RECT 137.145 123.335 137.315 123.505 ;
        RECT 137.605 123.335 137.775 123.505 ;
        RECT 138.065 123.335 138.235 123.505 ;
        RECT 138.525 123.335 138.695 123.505 ;
        RECT 138.985 123.335 139.155 123.505 ;
        RECT 50.665 120.615 50.835 120.785 ;
        RECT 51.125 120.615 51.295 120.785 ;
        RECT 51.585 120.615 51.755 120.785 ;
        RECT 52.045 120.615 52.215 120.785 ;
        RECT 52.505 120.615 52.675 120.785 ;
        RECT 52.965 120.615 53.135 120.785 ;
        RECT 53.425 120.615 53.595 120.785 ;
        RECT 53.885 120.615 54.055 120.785 ;
        RECT 54.345 120.615 54.515 120.785 ;
        RECT 54.805 120.615 54.975 120.785 ;
        RECT 55.265 120.615 55.435 120.785 ;
        RECT 55.725 120.615 55.895 120.785 ;
        RECT 56.185 120.615 56.355 120.785 ;
        RECT 56.645 120.615 56.815 120.785 ;
        RECT 57.105 120.615 57.275 120.785 ;
        RECT 57.565 120.615 57.735 120.785 ;
        RECT 58.025 120.615 58.195 120.785 ;
        RECT 58.485 120.615 58.655 120.785 ;
        RECT 58.945 120.615 59.115 120.785 ;
        RECT 59.405 120.615 59.575 120.785 ;
        RECT 59.865 120.615 60.035 120.785 ;
        RECT 60.325 120.615 60.495 120.785 ;
        RECT 60.785 120.615 60.955 120.785 ;
        RECT 61.245 120.615 61.415 120.785 ;
        RECT 61.705 120.615 61.875 120.785 ;
        RECT 62.165 120.615 62.335 120.785 ;
        RECT 62.625 120.615 62.795 120.785 ;
        RECT 63.085 120.615 63.255 120.785 ;
        RECT 63.545 120.615 63.715 120.785 ;
        RECT 64.005 120.615 64.175 120.785 ;
        RECT 64.465 120.615 64.635 120.785 ;
        RECT 64.925 120.615 65.095 120.785 ;
        RECT 65.385 120.615 65.555 120.785 ;
        RECT 65.845 120.615 66.015 120.785 ;
        RECT 66.305 120.615 66.475 120.785 ;
        RECT 66.765 120.615 66.935 120.785 ;
        RECT 67.225 120.615 67.395 120.785 ;
        RECT 67.685 120.615 67.855 120.785 ;
        RECT 68.145 120.615 68.315 120.785 ;
        RECT 68.605 120.615 68.775 120.785 ;
        RECT 69.065 120.615 69.235 120.785 ;
        RECT 69.525 120.615 69.695 120.785 ;
        RECT 69.985 120.615 70.155 120.785 ;
        RECT 70.445 120.615 70.615 120.785 ;
        RECT 70.905 120.615 71.075 120.785 ;
        RECT 71.365 120.615 71.535 120.785 ;
        RECT 71.825 120.615 71.995 120.785 ;
        RECT 72.285 120.615 72.455 120.785 ;
        RECT 72.745 120.615 72.915 120.785 ;
        RECT 73.205 120.615 73.375 120.785 ;
        RECT 73.665 120.615 73.835 120.785 ;
        RECT 74.125 120.615 74.295 120.785 ;
        RECT 74.585 120.615 74.755 120.785 ;
        RECT 75.045 120.615 75.215 120.785 ;
        RECT 75.505 120.615 75.675 120.785 ;
        RECT 75.965 120.615 76.135 120.785 ;
        RECT 76.425 120.615 76.595 120.785 ;
        RECT 76.885 120.615 77.055 120.785 ;
        RECT 77.345 120.615 77.515 120.785 ;
        RECT 77.805 120.615 77.975 120.785 ;
        RECT 78.265 120.615 78.435 120.785 ;
        RECT 78.725 120.615 78.895 120.785 ;
        RECT 79.185 120.615 79.355 120.785 ;
        RECT 79.645 120.615 79.815 120.785 ;
        RECT 80.105 120.615 80.275 120.785 ;
        RECT 80.565 120.615 80.735 120.785 ;
        RECT 81.025 120.615 81.195 120.785 ;
        RECT 81.485 120.615 81.655 120.785 ;
        RECT 81.945 120.615 82.115 120.785 ;
        RECT 82.405 120.615 82.575 120.785 ;
        RECT 82.865 120.615 83.035 120.785 ;
        RECT 83.325 120.615 83.495 120.785 ;
        RECT 83.785 120.615 83.955 120.785 ;
        RECT 84.245 120.615 84.415 120.785 ;
        RECT 84.705 120.615 84.875 120.785 ;
        RECT 85.165 120.615 85.335 120.785 ;
        RECT 85.625 120.615 85.795 120.785 ;
        RECT 86.085 120.615 86.255 120.785 ;
        RECT 86.545 120.615 86.715 120.785 ;
        RECT 87.005 120.615 87.175 120.785 ;
        RECT 87.465 120.615 87.635 120.785 ;
        RECT 87.925 120.615 88.095 120.785 ;
        RECT 88.385 120.615 88.555 120.785 ;
        RECT 88.845 120.615 89.015 120.785 ;
        RECT 89.305 120.615 89.475 120.785 ;
        RECT 89.765 120.615 89.935 120.785 ;
        RECT 90.225 120.615 90.395 120.785 ;
        RECT 90.685 120.615 90.855 120.785 ;
        RECT 91.145 120.615 91.315 120.785 ;
        RECT 91.605 120.615 91.775 120.785 ;
        RECT 92.065 120.615 92.235 120.785 ;
        RECT 92.525 120.615 92.695 120.785 ;
        RECT 92.985 120.615 93.155 120.785 ;
        RECT 93.445 120.615 93.615 120.785 ;
        RECT 93.905 120.615 94.075 120.785 ;
        RECT 94.365 120.615 94.535 120.785 ;
        RECT 94.825 120.615 94.995 120.785 ;
        RECT 95.285 120.615 95.455 120.785 ;
        RECT 95.745 120.615 95.915 120.785 ;
        RECT 96.205 120.615 96.375 120.785 ;
        RECT 96.665 120.615 96.835 120.785 ;
        RECT 97.125 120.615 97.295 120.785 ;
        RECT 97.585 120.615 97.755 120.785 ;
        RECT 98.045 120.615 98.215 120.785 ;
        RECT 98.505 120.615 98.675 120.785 ;
        RECT 98.965 120.615 99.135 120.785 ;
        RECT 99.425 120.615 99.595 120.785 ;
        RECT 99.885 120.615 100.055 120.785 ;
        RECT 100.345 120.615 100.515 120.785 ;
        RECT 100.805 120.615 100.975 120.785 ;
        RECT 101.265 120.615 101.435 120.785 ;
        RECT 101.725 120.615 101.895 120.785 ;
        RECT 102.185 120.615 102.355 120.785 ;
        RECT 102.645 120.615 102.815 120.785 ;
        RECT 103.105 120.615 103.275 120.785 ;
        RECT 103.565 120.615 103.735 120.785 ;
        RECT 104.025 120.615 104.195 120.785 ;
        RECT 104.485 120.615 104.655 120.785 ;
        RECT 104.945 120.615 105.115 120.785 ;
        RECT 105.405 120.615 105.575 120.785 ;
        RECT 105.865 120.615 106.035 120.785 ;
        RECT 106.325 120.615 106.495 120.785 ;
        RECT 106.785 120.615 106.955 120.785 ;
        RECT 107.245 120.615 107.415 120.785 ;
        RECT 107.705 120.615 107.875 120.785 ;
        RECT 108.165 120.615 108.335 120.785 ;
        RECT 108.625 120.615 108.795 120.785 ;
        RECT 109.085 120.615 109.255 120.785 ;
        RECT 109.545 120.615 109.715 120.785 ;
        RECT 110.005 120.615 110.175 120.785 ;
        RECT 110.465 120.615 110.635 120.785 ;
        RECT 110.925 120.615 111.095 120.785 ;
        RECT 111.385 120.615 111.555 120.785 ;
        RECT 111.845 120.615 112.015 120.785 ;
        RECT 112.305 120.615 112.475 120.785 ;
        RECT 112.765 120.615 112.935 120.785 ;
        RECT 113.225 120.615 113.395 120.785 ;
        RECT 113.685 120.615 113.855 120.785 ;
        RECT 114.145 120.615 114.315 120.785 ;
        RECT 114.605 120.615 114.775 120.785 ;
        RECT 115.065 120.615 115.235 120.785 ;
        RECT 115.525 120.615 115.695 120.785 ;
        RECT 115.985 120.615 116.155 120.785 ;
        RECT 116.445 120.615 116.615 120.785 ;
        RECT 116.905 120.615 117.075 120.785 ;
        RECT 117.365 120.615 117.535 120.785 ;
        RECT 117.825 120.615 117.995 120.785 ;
        RECT 118.285 120.615 118.455 120.785 ;
        RECT 118.745 120.615 118.915 120.785 ;
        RECT 119.205 120.615 119.375 120.785 ;
        RECT 119.665 120.615 119.835 120.785 ;
        RECT 120.125 120.615 120.295 120.785 ;
        RECT 120.585 120.615 120.755 120.785 ;
        RECT 121.045 120.615 121.215 120.785 ;
        RECT 121.505 120.615 121.675 120.785 ;
        RECT 121.965 120.615 122.135 120.785 ;
        RECT 122.425 120.615 122.595 120.785 ;
        RECT 122.885 120.615 123.055 120.785 ;
        RECT 123.345 120.615 123.515 120.785 ;
        RECT 123.805 120.615 123.975 120.785 ;
        RECT 124.265 120.615 124.435 120.785 ;
        RECT 124.725 120.615 124.895 120.785 ;
        RECT 125.185 120.615 125.355 120.785 ;
        RECT 125.645 120.615 125.815 120.785 ;
        RECT 126.105 120.615 126.275 120.785 ;
        RECT 126.565 120.615 126.735 120.785 ;
        RECT 127.025 120.615 127.195 120.785 ;
        RECT 127.485 120.615 127.655 120.785 ;
        RECT 127.945 120.615 128.115 120.785 ;
        RECT 128.405 120.615 128.575 120.785 ;
        RECT 128.865 120.615 129.035 120.785 ;
        RECT 129.325 120.615 129.495 120.785 ;
        RECT 129.785 120.615 129.955 120.785 ;
        RECT 130.245 120.615 130.415 120.785 ;
        RECT 130.705 120.615 130.875 120.785 ;
        RECT 131.165 120.615 131.335 120.785 ;
        RECT 131.625 120.615 131.795 120.785 ;
        RECT 132.085 120.615 132.255 120.785 ;
        RECT 132.545 120.615 132.715 120.785 ;
        RECT 133.005 120.615 133.175 120.785 ;
        RECT 133.465 120.615 133.635 120.785 ;
        RECT 133.925 120.615 134.095 120.785 ;
        RECT 134.385 120.615 134.555 120.785 ;
        RECT 134.845 120.615 135.015 120.785 ;
        RECT 135.305 120.615 135.475 120.785 ;
        RECT 135.765 120.615 135.935 120.785 ;
        RECT 136.225 120.615 136.395 120.785 ;
        RECT 136.685 120.615 136.855 120.785 ;
        RECT 137.145 120.615 137.315 120.785 ;
        RECT 137.605 120.615 137.775 120.785 ;
        RECT 138.065 120.615 138.235 120.785 ;
        RECT 138.525 120.615 138.695 120.785 ;
        RECT 138.985 120.615 139.155 120.785 ;
        RECT 50.665 117.895 50.835 118.065 ;
        RECT 51.125 117.895 51.295 118.065 ;
        RECT 51.585 117.895 51.755 118.065 ;
        RECT 52.045 117.895 52.215 118.065 ;
        RECT 52.505 117.895 52.675 118.065 ;
        RECT 52.965 117.895 53.135 118.065 ;
        RECT 53.425 117.895 53.595 118.065 ;
        RECT 53.885 117.895 54.055 118.065 ;
        RECT 54.345 117.895 54.515 118.065 ;
        RECT 54.805 117.895 54.975 118.065 ;
        RECT 55.265 117.895 55.435 118.065 ;
        RECT 55.725 117.895 55.895 118.065 ;
        RECT 56.185 117.895 56.355 118.065 ;
        RECT 56.645 117.895 56.815 118.065 ;
        RECT 57.105 117.895 57.275 118.065 ;
        RECT 57.565 117.895 57.735 118.065 ;
        RECT 58.025 117.895 58.195 118.065 ;
        RECT 58.485 117.895 58.655 118.065 ;
        RECT 58.945 117.895 59.115 118.065 ;
        RECT 59.405 117.895 59.575 118.065 ;
        RECT 59.865 117.895 60.035 118.065 ;
        RECT 60.325 117.895 60.495 118.065 ;
        RECT 60.785 117.895 60.955 118.065 ;
        RECT 61.245 117.895 61.415 118.065 ;
        RECT 61.705 117.895 61.875 118.065 ;
        RECT 62.165 117.895 62.335 118.065 ;
        RECT 62.625 117.895 62.795 118.065 ;
        RECT 63.085 117.895 63.255 118.065 ;
        RECT 63.545 117.895 63.715 118.065 ;
        RECT 64.005 117.895 64.175 118.065 ;
        RECT 64.465 117.895 64.635 118.065 ;
        RECT 64.925 117.895 65.095 118.065 ;
        RECT 65.385 117.895 65.555 118.065 ;
        RECT 65.845 117.895 66.015 118.065 ;
        RECT 66.305 117.895 66.475 118.065 ;
        RECT 66.765 117.895 66.935 118.065 ;
        RECT 67.225 117.895 67.395 118.065 ;
        RECT 67.685 117.895 67.855 118.065 ;
        RECT 68.145 117.895 68.315 118.065 ;
        RECT 68.605 117.895 68.775 118.065 ;
        RECT 69.065 117.895 69.235 118.065 ;
        RECT 69.525 117.895 69.695 118.065 ;
        RECT 69.985 117.895 70.155 118.065 ;
        RECT 70.445 117.895 70.615 118.065 ;
        RECT 70.905 117.895 71.075 118.065 ;
        RECT 71.365 117.895 71.535 118.065 ;
        RECT 71.825 117.895 71.995 118.065 ;
        RECT 72.285 117.895 72.455 118.065 ;
        RECT 72.745 117.895 72.915 118.065 ;
        RECT 73.205 117.895 73.375 118.065 ;
        RECT 73.665 117.895 73.835 118.065 ;
        RECT 74.125 117.895 74.295 118.065 ;
        RECT 74.585 117.895 74.755 118.065 ;
        RECT 75.045 117.895 75.215 118.065 ;
        RECT 75.505 117.895 75.675 118.065 ;
        RECT 75.965 117.895 76.135 118.065 ;
        RECT 76.425 117.895 76.595 118.065 ;
        RECT 76.885 117.895 77.055 118.065 ;
        RECT 77.345 117.895 77.515 118.065 ;
        RECT 77.805 117.895 77.975 118.065 ;
        RECT 78.265 117.895 78.435 118.065 ;
        RECT 78.725 117.895 78.895 118.065 ;
        RECT 79.185 117.895 79.355 118.065 ;
        RECT 79.645 117.895 79.815 118.065 ;
        RECT 80.105 117.895 80.275 118.065 ;
        RECT 80.565 117.895 80.735 118.065 ;
        RECT 81.025 117.895 81.195 118.065 ;
        RECT 81.485 117.895 81.655 118.065 ;
        RECT 81.945 117.895 82.115 118.065 ;
        RECT 82.405 117.895 82.575 118.065 ;
        RECT 82.865 117.895 83.035 118.065 ;
        RECT 83.325 117.895 83.495 118.065 ;
        RECT 83.785 117.895 83.955 118.065 ;
        RECT 84.245 117.895 84.415 118.065 ;
        RECT 84.705 117.895 84.875 118.065 ;
        RECT 85.165 117.895 85.335 118.065 ;
        RECT 85.625 117.895 85.795 118.065 ;
        RECT 86.085 117.895 86.255 118.065 ;
        RECT 86.545 117.895 86.715 118.065 ;
        RECT 87.005 117.895 87.175 118.065 ;
        RECT 87.465 117.895 87.635 118.065 ;
        RECT 87.925 117.895 88.095 118.065 ;
        RECT 88.385 117.895 88.555 118.065 ;
        RECT 88.845 117.895 89.015 118.065 ;
        RECT 89.305 117.895 89.475 118.065 ;
        RECT 89.765 117.895 89.935 118.065 ;
        RECT 90.225 117.895 90.395 118.065 ;
        RECT 90.685 117.895 90.855 118.065 ;
        RECT 91.145 117.895 91.315 118.065 ;
        RECT 91.605 117.895 91.775 118.065 ;
        RECT 92.065 117.895 92.235 118.065 ;
        RECT 92.525 117.895 92.695 118.065 ;
        RECT 92.985 117.895 93.155 118.065 ;
        RECT 93.445 117.895 93.615 118.065 ;
        RECT 93.905 117.895 94.075 118.065 ;
        RECT 94.365 117.895 94.535 118.065 ;
        RECT 94.825 117.895 94.995 118.065 ;
        RECT 95.285 117.895 95.455 118.065 ;
        RECT 95.745 117.895 95.915 118.065 ;
        RECT 96.205 117.895 96.375 118.065 ;
        RECT 96.665 117.895 96.835 118.065 ;
        RECT 97.125 117.895 97.295 118.065 ;
        RECT 97.585 117.895 97.755 118.065 ;
        RECT 98.045 117.895 98.215 118.065 ;
        RECT 98.505 117.895 98.675 118.065 ;
        RECT 98.965 117.895 99.135 118.065 ;
        RECT 99.425 117.895 99.595 118.065 ;
        RECT 99.885 117.895 100.055 118.065 ;
        RECT 100.345 117.895 100.515 118.065 ;
        RECT 100.805 117.895 100.975 118.065 ;
        RECT 101.265 117.895 101.435 118.065 ;
        RECT 101.725 117.895 101.895 118.065 ;
        RECT 102.185 117.895 102.355 118.065 ;
        RECT 102.645 117.895 102.815 118.065 ;
        RECT 103.105 117.895 103.275 118.065 ;
        RECT 103.565 117.895 103.735 118.065 ;
        RECT 104.025 117.895 104.195 118.065 ;
        RECT 104.485 117.895 104.655 118.065 ;
        RECT 104.945 117.895 105.115 118.065 ;
        RECT 105.405 117.895 105.575 118.065 ;
        RECT 105.865 117.895 106.035 118.065 ;
        RECT 106.325 117.895 106.495 118.065 ;
        RECT 106.785 117.895 106.955 118.065 ;
        RECT 107.245 117.895 107.415 118.065 ;
        RECT 107.705 117.895 107.875 118.065 ;
        RECT 108.165 117.895 108.335 118.065 ;
        RECT 108.625 117.895 108.795 118.065 ;
        RECT 109.085 117.895 109.255 118.065 ;
        RECT 109.545 117.895 109.715 118.065 ;
        RECT 110.005 117.895 110.175 118.065 ;
        RECT 110.465 117.895 110.635 118.065 ;
        RECT 110.925 117.895 111.095 118.065 ;
        RECT 111.385 117.895 111.555 118.065 ;
        RECT 111.845 117.895 112.015 118.065 ;
        RECT 112.305 117.895 112.475 118.065 ;
        RECT 112.765 117.895 112.935 118.065 ;
        RECT 113.225 117.895 113.395 118.065 ;
        RECT 113.685 117.895 113.855 118.065 ;
        RECT 114.145 117.895 114.315 118.065 ;
        RECT 114.605 117.895 114.775 118.065 ;
        RECT 115.065 117.895 115.235 118.065 ;
        RECT 115.525 117.895 115.695 118.065 ;
        RECT 115.985 117.895 116.155 118.065 ;
        RECT 116.445 117.895 116.615 118.065 ;
        RECT 116.905 117.895 117.075 118.065 ;
        RECT 117.365 117.895 117.535 118.065 ;
        RECT 117.825 117.895 117.995 118.065 ;
        RECT 118.285 117.895 118.455 118.065 ;
        RECT 118.745 117.895 118.915 118.065 ;
        RECT 119.205 117.895 119.375 118.065 ;
        RECT 119.665 117.895 119.835 118.065 ;
        RECT 120.125 117.895 120.295 118.065 ;
        RECT 120.585 117.895 120.755 118.065 ;
        RECT 121.045 117.895 121.215 118.065 ;
        RECT 121.505 117.895 121.675 118.065 ;
        RECT 121.965 117.895 122.135 118.065 ;
        RECT 122.425 117.895 122.595 118.065 ;
        RECT 122.885 117.895 123.055 118.065 ;
        RECT 123.345 117.895 123.515 118.065 ;
        RECT 123.805 117.895 123.975 118.065 ;
        RECT 124.265 117.895 124.435 118.065 ;
        RECT 124.725 117.895 124.895 118.065 ;
        RECT 125.185 117.895 125.355 118.065 ;
        RECT 125.645 117.895 125.815 118.065 ;
        RECT 126.105 117.895 126.275 118.065 ;
        RECT 126.565 117.895 126.735 118.065 ;
        RECT 127.025 117.895 127.195 118.065 ;
        RECT 127.485 117.895 127.655 118.065 ;
        RECT 127.945 117.895 128.115 118.065 ;
        RECT 128.405 117.895 128.575 118.065 ;
        RECT 128.865 117.895 129.035 118.065 ;
        RECT 129.325 117.895 129.495 118.065 ;
        RECT 129.785 117.895 129.955 118.065 ;
        RECT 130.245 117.895 130.415 118.065 ;
        RECT 130.705 117.895 130.875 118.065 ;
        RECT 131.165 117.895 131.335 118.065 ;
        RECT 131.625 117.895 131.795 118.065 ;
        RECT 132.085 117.895 132.255 118.065 ;
        RECT 132.545 117.895 132.715 118.065 ;
        RECT 133.005 117.895 133.175 118.065 ;
        RECT 133.465 117.895 133.635 118.065 ;
        RECT 133.925 117.895 134.095 118.065 ;
        RECT 134.385 117.895 134.555 118.065 ;
        RECT 134.845 117.895 135.015 118.065 ;
        RECT 135.305 117.895 135.475 118.065 ;
        RECT 135.765 117.895 135.935 118.065 ;
        RECT 136.225 117.895 136.395 118.065 ;
        RECT 136.685 117.895 136.855 118.065 ;
        RECT 137.145 117.895 137.315 118.065 ;
        RECT 137.605 117.895 137.775 118.065 ;
        RECT 138.065 117.895 138.235 118.065 ;
        RECT 138.525 117.895 138.695 118.065 ;
        RECT 138.985 117.895 139.155 118.065 ;
        RECT 50.665 115.175 50.835 115.345 ;
        RECT 51.125 115.175 51.295 115.345 ;
        RECT 51.585 115.175 51.755 115.345 ;
        RECT 52.045 115.175 52.215 115.345 ;
        RECT 52.505 115.175 52.675 115.345 ;
        RECT 52.965 115.175 53.135 115.345 ;
        RECT 53.425 115.175 53.595 115.345 ;
        RECT 53.885 115.175 54.055 115.345 ;
        RECT 54.345 115.175 54.515 115.345 ;
        RECT 54.805 115.175 54.975 115.345 ;
        RECT 55.265 115.175 55.435 115.345 ;
        RECT 55.725 115.175 55.895 115.345 ;
        RECT 56.185 115.175 56.355 115.345 ;
        RECT 56.645 115.175 56.815 115.345 ;
        RECT 57.105 115.175 57.275 115.345 ;
        RECT 57.565 115.175 57.735 115.345 ;
        RECT 58.025 115.175 58.195 115.345 ;
        RECT 58.485 115.175 58.655 115.345 ;
        RECT 58.945 115.175 59.115 115.345 ;
        RECT 59.405 115.175 59.575 115.345 ;
        RECT 59.865 115.175 60.035 115.345 ;
        RECT 60.325 115.175 60.495 115.345 ;
        RECT 60.785 115.175 60.955 115.345 ;
        RECT 61.245 115.175 61.415 115.345 ;
        RECT 61.705 115.175 61.875 115.345 ;
        RECT 62.165 115.175 62.335 115.345 ;
        RECT 62.625 115.175 62.795 115.345 ;
        RECT 63.085 115.175 63.255 115.345 ;
        RECT 63.545 115.175 63.715 115.345 ;
        RECT 64.005 115.175 64.175 115.345 ;
        RECT 64.465 115.175 64.635 115.345 ;
        RECT 64.925 115.175 65.095 115.345 ;
        RECT 65.385 115.175 65.555 115.345 ;
        RECT 65.845 115.175 66.015 115.345 ;
        RECT 66.305 115.175 66.475 115.345 ;
        RECT 66.765 115.175 66.935 115.345 ;
        RECT 67.225 115.175 67.395 115.345 ;
        RECT 67.685 115.175 67.855 115.345 ;
        RECT 68.145 115.175 68.315 115.345 ;
        RECT 68.605 115.175 68.775 115.345 ;
        RECT 69.065 115.175 69.235 115.345 ;
        RECT 69.525 115.175 69.695 115.345 ;
        RECT 69.985 115.175 70.155 115.345 ;
        RECT 70.445 115.175 70.615 115.345 ;
        RECT 70.905 115.175 71.075 115.345 ;
        RECT 71.365 115.175 71.535 115.345 ;
        RECT 71.825 115.175 71.995 115.345 ;
        RECT 72.285 115.175 72.455 115.345 ;
        RECT 72.745 115.175 72.915 115.345 ;
        RECT 73.205 115.175 73.375 115.345 ;
        RECT 73.665 115.175 73.835 115.345 ;
        RECT 74.125 115.175 74.295 115.345 ;
        RECT 74.585 115.175 74.755 115.345 ;
        RECT 75.045 115.175 75.215 115.345 ;
        RECT 75.505 115.175 75.675 115.345 ;
        RECT 75.965 115.175 76.135 115.345 ;
        RECT 76.425 115.175 76.595 115.345 ;
        RECT 76.885 115.175 77.055 115.345 ;
        RECT 77.345 115.175 77.515 115.345 ;
        RECT 77.805 115.175 77.975 115.345 ;
        RECT 78.265 115.175 78.435 115.345 ;
        RECT 78.725 115.175 78.895 115.345 ;
        RECT 79.185 115.175 79.355 115.345 ;
        RECT 79.645 115.175 79.815 115.345 ;
        RECT 80.105 115.175 80.275 115.345 ;
        RECT 80.565 115.175 80.735 115.345 ;
        RECT 81.025 115.175 81.195 115.345 ;
        RECT 81.485 115.175 81.655 115.345 ;
        RECT 81.945 115.175 82.115 115.345 ;
        RECT 82.405 115.175 82.575 115.345 ;
        RECT 82.865 115.175 83.035 115.345 ;
        RECT 83.325 115.175 83.495 115.345 ;
        RECT 83.785 115.175 83.955 115.345 ;
        RECT 84.245 115.175 84.415 115.345 ;
        RECT 84.705 115.175 84.875 115.345 ;
        RECT 85.165 115.175 85.335 115.345 ;
        RECT 85.625 115.175 85.795 115.345 ;
        RECT 86.085 115.175 86.255 115.345 ;
        RECT 86.545 115.175 86.715 115.345 ;
        RECT 87.005 115.175 87.175 115.345 ;
        RECT 87.465 115.175 87.635 115.345 ;
        RECT 87.925 115.175 88.095 115.345 ;
        RECT 88.385 115.175 88.555 115.345 ;
        RECT 88.845 115.175 89.015 115.345 ;
        RECT 89.305 115.175 89.475 115.345 ;
        RECT 89.765 115.175 89.935 115.345 ;
        RECT 90.225 115.175 90.395 115.345 ;
        RECT 90.685 115.175 90.855 115.345 ;
        RECT 91.145 115.175 91.315 115.345 ;
        RECT 91.605 115.175 91.775 115.345 ;
        RECT 92.065 115.175 92.235 115.345 ;
        RECT 92.525 115.175 92.695 115.345 ;
        RECT 92.985 115.175 93.155 115.345 ;
        RECT 93.445 115.175 93.615 115.345 ;
        RECT 93.905 115.175 94.075 115.345 ;
        RECT 94.365 115.175 94.535 115.345 ;
        RECT 94.825 115.175 94.995 115.345 ;
        RECT 95.285 115.175 95.455 115.345 ;
        RECT 95.745 115.175 95.915 115.345 ;
        RECT 96.205 115.175 96.375 115.345 ;
        RECT 96.665 115.175 96.835 115.345 ;
        RECT 97.125 115.175 97.295 115.345 ;
        RECT 97.585 115.175 97.755 115.345 ;
        RECT 98.045 115.175 98.215 115.345 ;
        RECT 98.505 115.175 98.675 115.345 ;
        RECT 98.965 115.175 99.135 115.345 ;
        RECT 99.425 115.175 99.595 115.345 ;
        RECT 99.885 115.175 100.055 115.345 ;
        RECT 100.345 115.175 100.515 115.345 ;
        RECT 100.805 115.175 100.975 115.345 ;
        RECT 101.265 115.175 101.435 115.345 ;
        RECT 101.725 115.175 101.895 115.345 ;
        RECT 102.185 115.175 102.355 115.345 ;
        RECT 102.645 115.175 102.815 115.345 ;
        RECT 103.105 115.175 103.275 115.345 ;
        RECT 103.565 115.175 103.735 115.345 ;
        RECT 104.025 115.175 104.195 115.345 ;
        RECT 104.485 115.175 104.655 115.345 ;
        RECT 104.945 115.175 105.115 115.345 ;
        RECT 105.405 115.175 105.575 115.345 ;
        RECT 105.865 115.175 106.035 115.345 ;
        RECT 106.325 115.175 106.495 115.345 ;
        RECT 106.785 115.175 106.955 115.345 ;
        RECT 107.245 115.175 107.415 115.345 ;
        RECT 107.705 115.175 107.875 115.345 ;
        RECT 108.165 115.175 108.335 115.345 ;
        RECT 108.625 115.175 108.795 115.345 ;
        RECT 109.085 115.175 109.255 115.345 ;
        RECT 109.545 115.175 109.715 115.345 ;
        RECT 110.005 115.175 110.175 115.345 ;
        RECT 110.465 115.175 110.635 115.345 ;
        RECT 110.925 115.175 111.095 115.345 ;
        RECT 111.385 115.175 111.555 115.345 ;
        RECT 111.845 115.175 112.015 115.345 ;
        RECT 112.305 115.175 112.475 115.345 ;
        RECT 112.765 115.175 112.935 115.345 ;
        RECT 113.225 115.175 113.395 115.345 ;
        RECT 113.685 115.175 113.855 115.345 ;
        RECT 114.145 115.175 114.315 115.345 ;
        RECT 114.605 115.175 114.775 115.345 ;
        RECT 115.065 115.175 115.235 115.345 ;
        RECT 115.525 115.175 115.695 115.345 ;
        RECT 115.985 115.175 116.155 115.345 ;
        RECT 116.445 115.175 116.615 115.345 ;
        RECT 116.905 115.175 117.075 115.345 ;
        RECT 117.365 115.175 117.535 115.345 ;
        RECT 117.825 115.175 117.995 115.345 ;
        RECT 118.285 115.175 118.455 115.345 ;
        RECT 118.745 115.175 118.915 115.345 ;
        RECT 119.205 115.175 119.375 115.345 ;
        RECT 119.665 115.175 119.835 115.345 ;
        RECT 120.125 115.175 120.295 115.345 ;
        RECT 120.585 115.175 120.755 115.345 ;
        RECT 121.045 115.175 121.215 115.345 ;
        RECT 121.505 115.175 121.675 115.345 ;
        RECT 121.965 115.175 122.135 115.345 ;
        RECT 122.425 115.175 122.595 115.345 ;
        RECT 122.885 115.175 123.055 115.345 ;
        RECT 123.345 115.175 123.515 115.345 ;
        RECT 123.805 115.175 123.975 115.345 ;
        RECT 124.265 115.175 124.435 115.345 ;
        RECT 124.725 115.175 124.895 115.345 ;
        RECT 125.185 115.175 125.355 115.345 ;
        RECT 125.645 115.175 125.815 115.345 ;
        RECT 126.105 115.175 126.275 115.345 ;
        RECT 126.565 115.175 126.735 115.345 ;
        RECT 127.025 115.175 127.195 115.345 ;
        RECT 127.485 115.175 127.655 115.345 ;
        RECT 127.945 115.175 128.115 115.345 ;
        RECT 128.405 115.175 128.575 115.345 ;
        RECT 128.865 115.175 129.035 115.345 ;
        RECT 129.325 115.175 129.495 115.345 ;
        RECT 129.785 115.175 129.955 115.345 ;
        RECT 130.245 115.175 130.415 115.345 ;
        RECT 130.705 115.175 130.875 115.345 ;
        RECT 131.165 115.175 131.335 115.345 ;
        RECT 131.625 115.175 131.795 115.345 ;
        RECT 132.085 115.175 132.255 115.345 ;
        RECT 132.545 115.175 132.715 115.345 ;
        RECT 133.005 115.175 133.175 115.345 ;
        RECT 133.465 115.175 133.635 115.345 ;
        RECT 133.925 115.175 134.095 115.345 ;
        RECT 134.385 115.175 134.555 115.345 ;
        RECT 134.845 115.175 135.015 115.345 ;
        RECT 135.305 115.175 135.475 115.345 ;
        RECT 135.765 115.175 135.935 115.345 ;
        RECT 136.225 115.175 136.395 115.345 ;
        RECT 136.685 115.175 136.855 115.345 ;
        RECT 137.145 115.175 137.315 115.345 ;
        RECT 137.605 115.175 137.775 115.345 ;
        RECT 138.065 115.175 138.235 115.345 ;
        RECT 138.525 115.175 138.695 115.345 ;
        RECT 138.985 115.175 139.155 115.345 ;
        RECT 50.665 112.455 50.835 112.625 ;
        RECT 51.125 112.455 51.295 112.625 ;
        RECT 51.585 112.455 51.755 112.625 ;
        RECT 52.045 112.455 52.215 112.625 ;
        RECT 52.505 112.455 52.675 112.625 ;
        RECT 52.965 112.455 53.135 112.625 ;
        RECT 53.425 112.455 53.595 112.625 ;
        RECT 53.885 112.455 54.055 112.625 ;
        RECT 54.345 112.455 54.515 112.625 ;
        RECT 54.805 112.455 54.975 112.625 ;
        RECT 55.265 112.455 55.435 112.625 ;
        RECT 55.725 112.455 55.895 112.625 ;
        RECT 56.185 112.455 56.355 112.625 ;
        RECT 56.645 112.455 56.815 112.625 ;
        RECT 57.105 112.455 57.275 112.625 ;
        RECT 57.565 112.455 57.735 112.625 ;
        RECT 58.025 112.455 58.195 112.625 ;
        RECT 58.485 112.455 58.655 112.625 ;
        RECT 58.945 112.455 59.115 112.625 ;
        RECT 59.405 112.455 59.575 112.625 ;
        RECT 59.865 112.455 60.035 112.625 ;
        RECT 60.325 112.455 60.495 112.625 ;
        RECT 60.785 112.455 60.955 112.625 ;
        RECT 61.245 112.455 61.415 112.625 ;
        RECT 61.705 112.455 61.875 112.625 ;
        RECT 62.165 112.455 62.335 112.625 ;
        RECT 62.625 112.455 62.795 112.625 ;
        RECT 63.085 112.455 63.255 112.625 ;
        RECT 63.545 112.455 63.715 112.625 ;
        RECT 64.005 112.455 64.175 112.625 ;
        RECT 64.465 112.455 64.635 112.625 ;
        RECT 64.925 112.455 65.095 112.625 ;
        RECT 65.385 112.455 65.555 112.625 ;
        RECT 65.845 112.455 66.015 112.625 ;
        RECT 66.305 112.455 66.475 112.625 ;
        RECT 66.765 112.455 66.935 112.625 ;
        RECT 67.225 112.455 67.395 112.625 ;
        RECT 67.685 112.455 67.855 112.625 ;
        RECT 68.145 112.455 68.315 112.625 ;
        RECT 68.605 112.455 68.775 112.625 ;
        RECT 69.065 112.455 69.235 112.625 ;
        RECT 69.525 112.455 69.695 112.625 ;
        RECT 69.985 112.455 70.155 112.625 ;
        RECT 70.445 112.455 70.615 112.625 ;
        RECT 70.905 112.455 71.075 112.625 ;
        RECT 71.365 112.455 71.535 112.625 ;
        RECT 71.825 112.455 71.995 112.625 ;
        RECT 72.285 112.455 72.455 112.625 ;
        RECT 72.745 112.455 72.915 112.625 ;
        RECT 73.205 112.455 73.375 112.625 ;
        RECT 73.665 112.455 73.835 112.625 ;
        RECT 74.125 112.455 74.295 112.625 ;
        RECT 74.585 112.455 74.755 112.625 ;
        RECT 75.045 112.455 75.215 112.625 ;
        RECT 75.505 112.455 75.675 112.625 ;
        RECT 75.965 112.455 76.135 112.625 ;
        RECT 76.425 112.455 76.595 112.625 ;
        RECT 76.885 112.455 77.055 112.625 ;
        RECT 77.345 112.455 77.515 112.625 ;
        RECT 77.805 112.455 77.975 112.625 ;
        RECT 78.265 112.455 78.435 112.625 ;
        RECT 78.725 112.455 78.895 112.625 ;
        RECT 79.185 112.455 79.355 112.625 ;
        RECT 79.645 112.455 79.815 112.625 ;
        RECT 80.105 112.455 80.275 112.625 ;
        RECT 80.565 112.455 80.735 112.625 ;
        RECT 81.025 112.455 81.195 112.625 ;
        RECT 81.485 112.455 81.655 112.625 ;
        RECT 81.945 112.455 82.115 112.625 ;
        RECT 82.405 112.455 82.575 112.625 ;
        RECT 82.865 112.455 83.035 112.625 ;
        RECT 83.325 112.455 83.495 112.625 ;
        RECT 83.785 112.455 83.955 112.625 ;
        RECT 84.245 112.455 84.415 112.625 ;
        RECT 84.705 112.455 84.875 112.625 ;
        RECT 85.165 112.455 85.335 112.625 ;
        RECT 85.625 112.455 85.795 112.625 ;
        RECT 86.085 112.455 86.255 112.625 ;
        RECT 86.545 112.455 86.715 112.625 ;
        RECT 87.005 112.455 87.175 112.625 ;
        RECT 87.465 112.455 87.635 112.625 ;
        RECT 87.925 112.455 88.095 112.625 ;
        RECT 88.385 112.455 88.555 112.625 ;
        RECT 88.845 112.455 89.015 112.625 ;
        RECT 89.305 112.455 89.475 112.625 ;
        RECT 89.765 112.455 89.935 112.625 ;
        RECT 90.225 112.455 90.395 112.625 ;
        RECT 90.685 112.455 90.855 112.625 ;
        RECT 91.145 112.455 91.315 112.625 ;
        RECT 91.605 112.455 91.775 112.625 ;
        RECT 92.065 112.455 92.235 112.625 ;
        RECT 92.525 112.455 92.695 112.625 ;
        RECT 92.985 112.455 93.155 112.625 ;
        RECT 93.445 112.455 93.615 112.625 ;
        RECT 93.905 112.455 94.075 112.625 ;
        RECT 94.365 112.455 94.535 112.625 ;
        RECT 94.825 112.455 94.995 112.625 ;
        RECT 95.285 112.455 95.455 112.625 ;
        RECT 95.745 112.455 95.915 112.625 ;
        RECT 96.205 112.455 96.375 112.625 ;
        RECT 96.665 112.455 96.835 112.625 ;
        RECT 97.125 112.455 97.295 112.625 ;
        RECT 97.585 112.455 97.755 112.625 ;
        RECT 98.045 112.455 98.215 112.625 ;
        RECT 98.505 112.455 98.675 112.625 ;
        RECT 98.965 112.455 99.135 112.625 ;
        RECT 99.425 112.455 99.595 112.625 ;
        RECT 99.885 112.455 100.055 112.625 ;
        RECT 100.345 112.455 100.515 112.625 ;
        RECT 100.805 112.455 100.975 112.625 ;
        RECT 101.265 112.455 101.435 112.625 ;
        RECT 101.725 112.455 101.895 112.625 ;
        RECT 102.185 112.455 102.355 112.625 ;
        RECT 102.645 112.455 102.815 112.625 ;
        RECT 103.105 112.455 103.275 112.625 ;
        RECT 103.565 112.455 103.735 112.625 ;
        RECT 104.025 112.455 104.195 112.625 ;
        RECT 104.485 112.455 104.655 112.625 ;
        RECT 104.945 112.455 105.115 112.625 ;
        RECT 105.405 112.455 105.575 112.625 ;
        RECT 105.865 112.455 106.035 112.625 ;
        RECT 106.325 112.455 106.495 112.625 ;
        RECT 106.785 112.455 106.955 112.625 ;
        RECT 107.245 112.455 107.415 112.625 ;
        RECT 107.705 112.455 107.875 112.625 ;
        RECT 108.165 112.455 108.335 112.625 ;
        RECT 108.625 112.455 108.795 112.625 ;
        RECT 109.085 112.455 109.255 112.625 ;
        RECT 109.545 112.455 109.715 112.625 ;
        RECT 110.005 112.455 110.175 112.625 ;
        RECT 110.465 112.455 110.635 112.625 ;
        RECT 110.925 112.455 111.095 112.625 ;
        RECT 111.385 112.455 111.555 112.625 ;
        RECT 111.845 112.455 112.015 112.625 ;
        RECT 112.305 112.455 112.475 112.625 ;
        RECT 112.765 112.455 112.935 112.625 ;
        RECT 113.225 112.455 113.395 112.625 ;
        RECT 113.685 112.455 113.855 112.625 ;
        RECT 114.145 112.455 114.315 112.625 ;
        RECT 114.605 112.455 114.775 112.625 ;
        RECT 115.065 112.455 115.235 112.625 ;
        RECT 115.525 112.455 115.695 112.625 ;
        RECT 115.985 112.455 116.155 112.625 ;
        RECT 116.445 112.455 116.615 112.625 ;
        RECT 116.905 112.455 117.075 112.625 ;
        RECT 117.365 112.455 117.535 112.625 ;
        RECT 117.825 112.455 117.995 112.625 ;
        RECT 118.285 112.455 118.455 112.625 ;
        RECT 118.745 112.455 118.915 112.625 ;
        RECT 119.205 112.455 119.375 112.625 ;
        RECT 119.665 112.455 119.835 112.625 ;
        RECT 120.125 112.455 120.295 112.625 ;
        RECT 120.585 112.455 120.755 112.625 ;
        RECT 121.045 112.455 121.215 112.625 ;
        RECT 121.505 112.455 121.675 112.625 ;
        RECT 121.965 112.455 122.135 112.625 ;
        RECT 122.425 112.455 122.595 112.625 ;
        RECT 122.885 112.455 123.055 112.625 ;
        RECT 123.345 112.455 123.515 112.625 ;
        RECT 123.805 112.455 123.975 112.625 ;
        RECT 124.265 112.455 124.435 112.625 ;
        RECT 124.725 112.455 124.895 112.625 ;
        RECT 125.185 112.455 125.355 112.625 ;
        RECT 125.645 112.455 125.815 112.625 ;
        RECT 126.105 112.455 126.275 112.625 ;
        RECT 126.565 112.455 126.735 112.625 ;
        RECT 127.025 112.455 127.195 112.625 ;
        RECT 127.485 112.455 127.655 112.625 ;
        RECT 127.945 112.455 128.115 112.625 ;
        RECT 128.405 112.455 128.575 112.625 ;
        RECT 128.865 112.455 129.035 112.625 ;
        RECT 129.325 112.455 129.495 112.625 ;
        RECT 129.785 112.455 129.955 112.625 ;
        RECT 130.245 112.455 130.415 112.625 ;
        RECT 130.705 112.455 130.875 112.625 ;
        RECT 131.165 112.455 131.335 112.625 ;
        RECT 131.625 112.455 131.795 112.625 ;
        RECT 132.085 112.455 132.255 112.625 ;
        RECT 132.545 112.455 132.715 112.625 ;
        RECT 133.005 112.455 133.175 112.625 ;
        RECT 133.465 112.455 133.635 112.625 ;
        RECT 133.925 112.455 134.095 112.625 ;
        RECT 134.385 112.455 134.555 112.625 ;
        RECT 134.845 112.455 135.015 112.625 ;
        RECT 135.305 112.455 135.475 112.625 ;
        RECT 135.765 112.455 135.935 112.625 ;
        RECT 136.225 112.455 136.395 112.625 ;
        RECT 136.685 112.455 136.855 112.625 ;
        RECT 137.145 112.455 137.315 112.625 ;
        RECT 137.605 112.455 137.775 112.625 ;
        RECT 138.065 112.455 138.235 112.625 ;
        RECT 138.525 112.455 138.695 112.625 ;
        RECT 138.985 112.455 139.155 112.625 ;
        RECT 50.665 109.735 50.835 109.905 ;
        RECT 51.125 109.735 51.295 109.905 ;
        RECT 51.585 109.735 51.755 109.905 ;
        RECT 52.045 109.735 52.215 109.905 ;
        RECT 52.505 109.735 52.675 109.905 ;
        RECT 52.965 109.735 53.135 109.905 ;
        RECT 53.425 109.735 53.595 109.905 ;
        RECT 53.885 109.735 54.055 109.905 ;
        RECT 54.345 109.735 54.515 109.905 ;
        RECT 54.805 109.735 54.975 109.905 ;
        RECT 55.265 109.735 55.435 109.905 ;
        RECT 55.725 109.735 55.895 109.905 ;
        RECT 56.185 109.735 56.355 109.905 ;
        RECT 56.645 109.735 56.815 109.905 ;
        RECT 57.105 109.735 57.275 109.905 ;
        RECT 57.565 109.735 57.735 109.905 ;
        RECT 58.025 109.735 58.195 109.905 ;
        RECT 58.485 109.735 58.655 109.905 ;
        RECT 58.945 109.735 59.115 109.905 ;
        RECT 59.405 109.735 59.575 109.905 ;
        RECT 59.865 109.735 60.035 109.905 ;
        RECT 60.325 109.735 60.495 109.905 ;
        RECT 60.785 109.735 60.955 109.905 ;
        RECT 61.245 109.735 61.415 109.905 ;
        RECT 61.705 109.735 61.875 109.905 ;
        RECT 62.165 109.735 62.335 109.905 ;
        RECT 62.625 109.735 62.795 109.905 ;
        RECT 63.085 109.735 63.255 109.905 ;
        RECT 63.545 109.735 63.715 109.905 ;
        RECT 64.005 109.735 64.175 109.905 ;
        RECT 64.465 109.735 64.635 109.905 ;
        RECT 64.925 109.735 65.095 109.905 ;
        RECT 65.385 109.735 65.555 109.905 ;
        RECT 65.845 109.735 66.015 109.905 ;
        RECT 66.305 109.735 66.475 109.905 ;
        RECT 66.765 109.735 66.935 109.905 ;
        RECT 67.225 109.735 67.395 109.905 ;
        RECT 67.685 109.735 67.855 109.905 ;
        RECT 68.145 109.735 68.315 109.905 ;
        RECT 68.605 109.735 68.775 109.905 ;
        RECT 69.065 109.735 69.235 109.905 ;
        RECT 69.525 109.735 69.695 109.905 ;
        RECT 69.985 109.735 70.155 109.905 ;
        RECT 70.445 109.735 70.615 109.905 ;
        RECT 70.905 109.735 71.075 109.905 ;
        RECT 71.365 109.735 71.535 109.905 ;
        RECT 71.825 109.735 71.995 109.905 ;
        RECT 72.285 109.735 72.455 109.905 ;
        RECT 72.745 109.735 72.915 109.905 ;
        RECT 73.205 109.735 73.375 109.905 ;
        RECT 73.665 109.735 73.835 109.905 ;
        RECT 74.125 109.735 74.295 109.905 ;
        RECT 74.585 109.735 74.755 109.905 ;
        RECT 75.045 109.735 75.215 109.905 ;
        RECT 75.505 109.735 75.675 109.905 ;
        RECT 75.965 109.735 76.135 109.905 ;
        RECT 76.425 109.735 76.595 109.905 ;
        RECT 76.885 109.735 77.055 109.905 ;
        RECT 77.345 109.735 77.515 109.905 ;
        RECT 77.805 109.735 77.975 109.905 ;
        RECT 78.265 109.735 78.435 109.905 ;
        RECT 78.725 109.735 78.895 109.905 ;
        RECT 79.185 109.735 79.355 109.905 ;
        RECT 79.645 109.735 79.815 109.905 ;
        RECT 80.105 109.735 80.275 109.905 ;
        RECT 80.565 109.735 80.735 109.905 ;
        RECT 81.025 109.735 81.195 109.905 ;
        RECT 81.485 109.735 81.655 109.905 ;
        RECT 81.945 109.735 82.115 109.905 ;
        RECT 82.405 109.735 82.575 109.905 ;
        RECT 82.865 109.735 83.035 109.905 ;
        RECT 83.325 109.735 83.495 109.905 ;
        RECT 83.785 109.735 83.955 109.905 ;
        RECT 84.245 109.735 84.415 109.905 ;
        RECT 84.705 109.735 84.875 109.905 ;
        RECT 85.165 109.735 85.335 109.905 ;
        RECT 85.625 109.735 85.795 109.905 ;
        RECT 86.085 109.735 86.255 109.905 ;
        RECT 86.545 109.735 86.715 109.905 ;
        RECT 87.005 109.735 87.175 109.905 ;
        RECT 87.465 109.735 87.635 109.905 ;
        RECT 87.925 109.735 88.095 109.905 ;
        RECT 88.385 109.735 88.555 109.905 ;
        RECT 88.845 109.735 89.015 109.905 ;
        RECT 89.305 109.735 89.475 109.905 ;
        RECT 89.765 109.735 89.935 109.905 ;
        RECT 90.225 109.735 90.395 109.905 ;
        RECT 90.685 109.735 90.855 109.905 ;
        RECT 91.145 109.735 91.315 109.905 ;
        RECT 91.605 109.735 91.775 109.905 ;
        RECT 92.065 109.735 92.235 109.905 ;
        RECT 92.525 109.735 92.695 109.905 ;
        RECT 92.985 109.735 93.155 109.905 ;
        RECT 93.445 109.735 93.615 109.905 ;
        RECT 93.905 109.735 94.075 109.905 ;
        RECT 94.365 109.735 94.535 109.905 ;
        RECT 94.825 109.735 94.995 109.905 ;
        RECT 95.285 109.735 95.455 109.905 ;
        RECT 95.745 109.735 95.915 109.905 ;
        RECT 96.205 109.735 96.375 109.905 ;
        RECT 96.665 109.735 96.835 109.905 ;
        RECT 97.125 109.735 97.295 109.905 ;
        RECT 97.585 109.735 97.755 109.905 ;
        RECT 98.045 109.735 98.215 109.905 ;
        RECT 98.505 109.735 98.675 109.905 ;
        RECT 98.965 109.735 99.135 109.905 ;
        RECT 99.425 109.735 99.595 109.905 ;
        RECT 99.885 109.735 100.055 109.905 ;
        RECT 100.345 109.735 100.515 109.905 ;
        RECT 100.805 109.735 100.975 109.905 ;
        RECT 101.265 109.735 101.435 109.905 ;
        RECT 101.725 109.735 101.895 109.905 ;
        RECT 102.185 109.735 102.355 109.905 ;
        RECT 102.645 109.735 102.815 109.905 ;
        RECT 103.105 109.735 103.275 109.905 ;
        RECT 103.565 109.735 103.735 109.905 ;
        RECT 104.025 109.735 104.195 109.905 ;
        RECT 104.485 109.735 104.655 109.905 ;
        RECT 104.945 109.735 105.115 109.905 ;
        RECT 105.405 109.735 105.575 109.905 ;
        RECT 105.865 109.735 106.035 109.905 ;
        RECT 106.325 109.735 106.495 109.905 ;
        RECT 106.785 109.735 106.955 109.905 ;
        RECT 107.245 109.735 107.415 109.905 ;
        RECT 107.705 109.735 107.875 109.905 ;
        RECT 108.165 109.735 108.335 109.905 ;
        RECT 108.625 109.735 108.795 109.905 ;
        RECT 109.085 109.735 109.255 109.905 ;
        RECT 109.545 109.735 109.715 109.905 ;
        RECT 110.005 109.735 110.175 109.905 ;
        RECT 110.465 109.735 110.635 109.905 ;
        RECT 110.925 109.735 111.095 109.905 ;
        RECT 111.385 109.735 111.555 109.905 ;
        RECT 111.845 109.735 112.015 109.905 ;
        RECT 112.305 109.735 112.475 109.905 ;
        RECT 112.765 109.735 112.935 109.905 ;
        RECT 113.225 109.735 113.395 109.905 ;
        RECT 113.685 109.735 113.855 109.905 ;
        RECT 114.145 109.735 114.315 109.905 ;
        RECT 114.605 109.735 114.775 109.905 ;
        RECT 115.065 109.735 115.235 109.905 ;
        RECT 115.525 109.735 115.695 109.905 ;
        RECT 115.985 109.735 116.155 109.905 ;
        RECT 116.445 109.735 116.615 109.905 ;
        RECT 116.905 109.735 117.075 109.905 ;
        RECT 117.365 109.735 117.535 109.905 ;
        RECT 117.825 109.735 117.995 109.905 ;
        RECT 118.285 109.735 118.455 109.905 ;
        RECT 118.745 109.735 118.915 109.905 ;
        RECT 119.205 109.735 119.375 109.905 ;
        RECT 119.665 109.735 119.835 109.905 ;
        RECT 120.125 109.735 120.295 109.905 ;
        RECT 120.585 109.735 120.755 109.905 ;
        RECT 121.045 109.735 121.215 109.905 ;
        RECT 121.505 109.735 121.675 109.905 ;
        RECT 121.965 109.735 122.135 109.905 ;
        RECT 122.425 109.735 122.595 109.905 ;
        RECT 122.885 109.735 123.055 109.905 ;
        RECT 123.345 109.735 123.515 109.905 ;
        RECT 123.805 109.735 123.975 109.905 ;
        RECT 124.265 109.735 124.435 109.905 ;
        RECT 124.725 109.735 124.895 109.905 ;
        RECT 125.185 109.735 125.355 109.905 ;
        RECT 125.645 109.735 125.815 109.905 ;
        RECT 126.105 109.735 126.275 109.905 ;
        RECT 126.565 109.735 126.735 109.905 ;
        RECT 127.025 109.735 127.195 109.905 ;
        RECT 127.485 109.735 127.655 109.905 ;
        RECT 127.945 109.735 128.115 109.905 ;
        RECT 128.405 109.735 128.575 109.905 ;
        RECT 128.865 109.735 129.035 109.905 ;
        RECT 129.325 109.735 129.495 109.905 ;
        RECT 129.785 109.735 129.955 109.905 ;
        RECT 130.245 109.735 130.415 109.905 ;
        RECT 130.705 109.735 130.875 109.905 ;
        RECT 131.165 109.735 131.335 109.905 ;
        RECT 131.625 109.735 131.795 109.905 ;
        RECT 132.085 109.735 132.255 109.905 ;
        RECT 132.545 109.735 132.715 109.905 ;
        RECT 133.005 109.735 133.175 109.905 ;
        RECT 133.465 109.735 133.635 109.905 ;
        RECT 133.925 109.735 134.095 109.905 ;
        RECT 134.385 109.735 134.555 109.905 ;
        RECT 134.845 109.735 135.015 109.905 ;
        RECT 135.305 109.735 135.475 109.905 ;
        RECT 135.765 109.735 135.935 109.905 ;
        RECT 136.225 109.735 136.395 109.905 ;
        RECT 136.685 109.735 136.855 109.905 ;
        RECT 137.145 109.735 137.315 109.905 ;
        RECT 137.605 109.735 137.775 109.905 ;
        RECT 138.065 109.735 138.235 109.905 ;
        RECT 138.525 109.735 138.695 109.905 ;
        RECT 138.985 109.735 139.155 109.905 ;
        RECT 65.385 108.545 65.555 108.715 ;
        RECT 65.845 108.545 66.015 108.715 ;
        RECT 66.765 108.545 66.935 108.715 ;
        RECT 50.665 107.015 50.835 107.185 ;
        RECT 51.125 107.015 51.295 107.185 ;
        RECT 51.585 107.015 51.755 107.185 ;
        RECT 52.045 107.015 52.215 107.185 ;
        RECT 52.505 107.015 52.675 107.185 ;
        RECT 52.965 107.015 53.135 107.185 ;
        RECT 53.425 107.015 53.595 107.185 ;
        RECT 53.885 107.015 54.055 107.185 ;
        RECT 54.345 107.015 54.515 107.185 ;
        RECT 54.805 107.015 54.975 107.185 ;
        RECT 55.265 107.015 55.435 107.185 ;
        RECT 55.725 107.015 55.895 107.185 ;
        RECT 56.185 107.015 56.355 107.185 ;
        RECT 56.645 107.015 56.815 107.185 ;
        RECT 57.105 107.015 57.275 107.185 ;
        RECT 57.565 107.015 57.735 107.185 ;
        RECT 58.025 107.015 58.195 107.185 ;
        RECT 58.485 107.015 58.655 107.185 ;
        RECT 58.945 107.015 59.115 107.185 ;
        RECT 59.405 107.015 59.575 107.185 ;
        RECT 59.865 107.015 60.035 107.185 ;
        RECT 60.325 107.015 60.495 107.185 ;
        RECT 60.785 107.015 60.955 107.185 ;
        RECT 61.245 107.015 61.415 107.185 ;
        RECT 61.705 107.015 61.875 107.185 ;
        RECT 62.165 107.015 62.335 107.185 ;
        RECT 62.625 107.015 62.795 107.185 ;
        RECT 63.085 107.015 63.255 107.185 ;
        RECT 63.545 107.015 63.715 107.185 ;
        RECT 64.005 107.015 64.175 107.185 ;
        RECT 64.465 107.015 64.635 107.185 ;
        RECT 64.925 107.015 65.095 107.185 ;
        RECT 65.385 107.015 65.555 107.185 ;
        RECT 65.845 107.015 66.015 107.185 ;
        RECT 66.305 107.015 66.475 107.185 ;
        RECT 66.765 107.015 66.935 107.185 ;
        RECT 67.225 107.015 67.395 107.185 ;
        RECT 67.685 107.015 67.855 107.185 ;
        RECT 68.145 107.015 68.315 107.185 ;
        RECT 68.605 107.015 68.775 107.185 ;
        RECT 69.065 107.015 69.235 107.185 ;
        RECT 69.525 107.015 69.695 107.185 ;
        RECT 69.985 107.015 70.155 107.185 ;
        RECT 70.445 107.015 70.615 107.185 ;
        RECT 70.905 107.015 71.075 107.185 ;
        RECT 71.365 107.015 71.535 107.185 ;
        RECT 71.825 107.015 71.995 107.185 ;
        RECT 72.285 107.015 72.455 107.185 ;
        RECT 72.745 107.015 72.915 107.185 ;
        RECT 73.205 107.015 73.375 107.185 ;
        RECT 73.665 107.015 73.835 107.185 ;
        RECT 74.125 107.015 74.295 107.185 ;
        RECT 74.585 107.015 74.755 107.185 ;
        RECT 75.045 107.015 75.215 107.185 ;
        RECT 75.505 107.015 75.675 107.185 ;
        RECT 75.965 107.015 76.135 107.185 ;
        RECT 76.425 107.015 76.595 107.185 ;
        RECT 76.885 107.015 77.055 107.185 ;
        RECT 77.345 107.015 77.515 107.185 ;
        RECT 77.805 107.015 77.975 107.185 ;
        RECT 78.265 107.015 78.435 107.185 ;
        RECT 78.725 107.015 78.895 107.185 ;
        RECT 79.185 107.015 79.355 107.185 ;
        RECT 79.645 107.015 79.815 107.185 ;
        RECT 80.105 107.015 80.275 107.185 ;
        RECT 80.565 107.015 80.735 107.185 ;
        RECT 81.025 107.015 81.195 107.185 ;
        RECT 81.485 107.015 81.655 107.185 ;
        RECT 81.945 107.015 82.115 107.185 ;
        RECT 82.405 107.015 82.575 107.185 ;
        RECT 82.865 107.015 83.035 107.185 ;
        RECT 83.325 107.015 83.495 107.185 ;
        RECT 83.785 107.015 83.955 107.185 ;
        RECT 84.245 107.015 84.415 107.185 ;
        RECT 84.705 107.015 84.875 107.185 ;
        RECT 85.165 107.015 85.335 107.185 ;
        RECT 85.625 107.015 85.795 107.185 ;
        RECT 86.085 107.015 86.255 107.185 ;
        RECT 86.545 107.015 86.715 107.185 ;
        RECT 87.005 107.015 87.175 107.185 ;
        RECT 87.465 107.015 87.635 107.185 ;
        RECT 87.925 107.015 88.095 107.185 ;
        RECT 88.385 107.015 88.555 107.185 ;
        RECT 88.845 107.015 89.015 107.185 ;
        RECT 89.305 107.015 89.475 107.185 ;
        RECT 89.765 107.015 89.935 107.185 ;
        RECT 90.225 107.015 90.395 107.185 ;
        RECT 90.685 107.015 90.855 107.185 ;
        RECT 91.145 107.015 91.315 107.185 ;
        RECT 91.605 107.015 91.775 107.185 ;
        RECT 92.065 107.015 92.235 107.185 ;
        RECT 92.525 107.015 92.695 107.185 ;
        RECT 92.985 107.015 93.155 107.185 ;
        RECT 93.445 107.015 93.615 107.185 ;
        RECT 93.905 107.015 94.075 107.185 ;
        RECT 94.365 107.015 94.535 107.185 ;
        RECT 94.825 107.015 94.995 107.185 ;
        RECT 95.285 107.015 95.455 107.185 ;
        RECT 95.745 107.015 95.915 107.185 ;
        RECT 96.205 107.015 96.375 107.185 ;
        RECT 96.665 107.015 96.835 107.185 ;
        RECT 97.125 107.015 97.295 107.185 ;
        RECT 97.585 107.015 97.755 107.185 ;
        RECT 98.045 107.015 98.215 107.185 ;
        RECT 98.505 107.015 98.675 107.185 ;
        RECT 98.965 107.015 99.135 107.185 ;
        RECT 99.425 107.015 99.595 107.185 ;
        RECT 99.885 107.015 100.055 107.185 ;
        RECT 100.345 107.015 100.515 107.185 ;
        RECT 100.805 107.015 100.975 107.185 ;
        RECT 101.265 107.015 101.435 107.185 ;
        RECT 101.725 107.015 101.895 107.185 ;
        RECT 102.185 107.015 102.355 107.185 ;
        RECT 102.645 107.015 102.815 107.185 ;
        RECT 103.105 107.015 103.275 107.185 ;
        RECT 103.565 107.015 103.735 107.185 ;
        RECT 104.025 107.015 104.195 107.185 ;
        RECT 104.485 107.015 104.655 107.185 ;
        RECT 104.945 107.015 105.115 107.185 ;
        RECT 105.405 107.015 105.575 107.185 ;
        RECT 105.865 107.015 106.035 107.185 ;
        RECT 106.325 107.015 106.495 107.185 ;
        RECT 106.785 107.015 106.955 107.185 ;
        RECT 107.245 107.015 107.415 107.185 ;
        RECT 107.705 107.015 107.875 107.185 ;
        RECT 108.165 107.015 108.335 107.185 ;
        RECT 108.625 107.015 108.795 107.185 ;
        RECT 109.085 107.015 109.255 107.185 ;
        RECT 109.545 107.015 109.715 107.185 ;
        RECT 110.005 107.015 110.175 107.185 ;
        RECT 110.465 107.015 110.635 107.185 ;
        RECT 110.925 107.015 111.095 107.185 ;
        RECT 111.385 107.015 111.555 107.185 ;
        RECT 111.845 107.015 112.015 107.185 ;
        RECT 112.305 107.015 112.475 107.185 ;
        RECT 112.765 107.015 112.935 107.185 ;
        RECT 113.225 107.015 113.395 107.185 ;
        RECT 113.685 107.015 113.855 107.185 ;
        RECT 114.145 107.015 114.315 107.185 ;
        RECT 114.605 107.015 114.775 107.185 ;
        RECT 115.065 107.015 115.235 107.185 ;
        RECT 115.525 107.015 115.695 107.185 ;
        RECT 115.985 107.015 116.155 107.185 ;
        RECT 116.445 107.015 116.615 107.185 ;
        RECT 116.905 107.015 117.075 107.185 ;
        RECT 117.365 107.015 117.535 107.185 ;
        RECT 117.825 107.015 117.995 107.185 ;
        RECT 118.285 107.015 118.455 107.185 ;
        RECT 118.745 107.015 118.915 107.185 ;
        RECT 119.205 107.015 119.375 107.185 ;
        RECT 119.665 107.015 119.835 107.185 ;
        RECT 120.125 107.015 120.295 107.185 ;
        RECT 120.585 107.015 120.755 107.185 ;
        RECT 121.045 107.015 121.215 107.185 ;
        RECT 121.505 107.015 121.675 107.185 ;
        RECT 121.965 107.015 122.135 107.185 ;
        RECT 122.425 107.015 122.595 107.185 ;
        RECT 122.885 107.015 123.055 107.185 ;
        RECT 123.345 107.015 123.515 107.185 ;
        RECT 123.805 107.015 123.975 107.185 ;
        RECT 124.265 107.015 124.435 107.185 ;
        RECT 124.725 107.015 124.895 107.185 ;
        RECT 125.185 107.015 125.355 107.185 ;
        RECT 125.645 107.015 125.815 107.185 ;
        RECT 126.105 107.015 126.275 107.185 ;
        RECT 126.565 107.015 126.735 107.185 ;
        RECT 127.025 107.015 127.195 107.185 ;
        RECT 127.485 107.015 127.655 107.185 ;
        RECT 127.945 107.015 128.115 107.185 ;
        RECT 128.405 107.015 128.575 107.185 ;
        RECT 128.865 107.015 129.035 107.185 ;
        RECT 129.325 107.015 129.495 107.185 ;
        RECT 129.785 107.015 129.955 107.185 ;
        RECT 130.245 107.015 130.415 107.185 ;
        RECT 130.705 107.015 130.875 107.185 ;
        RECT 131.165 107.015 131.335 107.185 ;
        RECT 131.625 107.015 131.795 107.185 ;
        RECT 132.085 107.015 132.255 107.185 ;
        RECT 132.545 107.015 132.715 107.185 ;
        RECT 133.005 107.015 133.175 107.185 ;
        RECT 133.465 107.015 133.635 107.185 ;
        RECT 133.925 107.015 134.095 107.185 ;
        RECT 134.385 107.015 134.555 107.185 ;
        RECT 134.845 107.015 135.015 107.185 ;
        RECT 135.305 107.015 135.475 107.185 ;
        RECT 135.765 107.015 135.935 107.185 ;
        RECT 136.225 107.015 136.395 107.185 ;
        RECT 136.685 107.015 136.855 107.185 ;
        RECT 137.145 107.015 137.315 107.185 ;
        RECT 137.605 107.015 137.775 107.185 ;
        RECT 138.065 107.015 138.235 107.185 ;
        RECT 138.525 107.015 138.695 107.185 ;
        RECT 138.985 107.015 139.155 107.185 ;
        RECT 58.025 105.825 58.195 105.995 ;
        RECT 57.105 105.485 57.275 105.655 ;
        RECT 57.565 105.485 57.735 105.655 ;
        RECT 58.485 105.485 58.655 105.655 ;
        RECT 61.245 105.825 61.415 105.995 ;
        RECT 58.945 105.145 59.115 105.315 ;
        RECT 62.165 105.485 62.335 105.655 ;
        RECT 50.665 104.295 50.835 104.465 ;
        RECT 51.125 104.295 51.295 104.465 ;
        RECT 51.585 104.295 51.755 104.465 ;
        RECT 52.045 104.295 52.215 104.465 ;
        RECT 52.505 104.295 52.675 104.465 ;
        RECT 52.965 104.295 53.135 104.465 ;
        RECT 53.425 104.295 53.595 104.465 ;
        RECT 53.885 104.295 54.055 104.465 ;
        RECT 54.345 104.295 54.515 104.465 ;
        RECT 54.805 104.295 54.975 104.465 ;
        RECT 55.265 104.295 55.435 104.465 ;
        RECT 55.725 104.295 55.895 104.465 ;
        RECT 56.185 104.295 56.355 104.465 ;
        RECT 56.645 104.295 56.815 104.465 ;
        RECT 57.105 104.295 57.275 104.465 ;
        RECT 57.565 104.295 57.735 104.465 ;
        RECT 58.025 104.295 58.195 104.465 ;
        RECT 58.485 104.295 58.655 104.465 ;
        RECT 58.945 104.295 59.115 104.465 ;
        RECT 59.405 104.295 59.575 104.465 ;
        RECT 59.865 104.295 60.035 104.465 ;
        RECT 60.325 104.295 60.495 104.465 ;
        RECT 60.785 104.295 60.955 104.465 ;
        RECT 61.245 104.295 61.415 104.465 ;
        RECT 61.705 104.295 61.875 104.465 ;
        RECT 62.165 104.295 62.335 104.465 ;
        RECT 62.625 104.295 62.795 104.465 ;
        RECT 63.085 104.295 63.255 104.465 ;
        RECT 63.545 104.295 63.715 104.465 ;
        RECT 64.005 104.295 64.175 104.465 ;
        RECT 64.465 104.295 64.635 104.465 ;
        RECT 64.925 104.295 65.095 104.465 ;
        RECT 65.385 104.295 65.555 104.465 ;
        RECT 65.845 104.295 66.015 104.465 ;
        RECT 66.305 104.295 66.475 104.465 ;
        RECT 66.765 104.295 66.935 104.465 ;
        RECT 67.225 104.295 67.395 104.465 ;
        RECT 67.685 104.295 67.855 104.465 ;
        RECT 68.145 104.295 68.315 104.465 ;
        RECT 68.605 104.295 68.775 104.465 ;
        RECT 69.065 104.295 69.235 104.465 ;
        RECT 69.525 104.295 69.695 104.465 ;
        RECT 69.985 104.295 70.155 104.465 ;
        RECT 70.445 104.295 70.615 104.465 ;
        RECT 70.905 104.295 71.075 104.465 ;
        RECT 71.365 104.295 71.535 104.465 ;
        RECT 71.825 104.295 71.995 104.465 ;
        RECT 72.285 104.295 72.455 104.465 ;
        RECT 72.745 104.295 72.915 104.465 ;
        RECT 73.205 104.295 73.375 104.465 ;
        RECT 73.665 104.295 73.835 104.465 ;
        RECT 74.125 104.295 74.295 104.465 ;
        RECT 74.585 104.295 74.755 104.465 ;
        RECT 75.045 104.295 75.215 104.465 ;
        RECT 75.505 104.295 75.675 104.465 ;
        RECT 75.965 104.295 76.135 104.465 ;
        RECT 76.425 104.295 76.595 104.465 ;
        RECT 76.885 104.295 77.055 104.465 ;
        RECT 77.345 104.295 77.515 104.465 ;
        RECT 77.805 104.295 77.975 104.465 ;
        RECT 78.265 104.295 78.435 104.465 ;
        RECT 78.725 104.295 78.895 104.465 ;
        RECT 79.185 104.295 79.355 104.465 ;
        RECT 79.645 104.295 79.815 104.465 ;
        RECT 80.105 104.295 80.275 104.465 ;
        RECT 80.565 104.295 80.735 104.465 ;
        RECT 81.025 104.295 81.195 104.465 ;
        RECT 81.485 104.295 81.655 104.465 ;
        RECT 81.945 104.295 82.115 104.465 ;
        RECT 82.405 104.295 82.575 104.465 ;
        RECT 82.865 104.295 83.035 104.465 ;
        RECT 83.325 104.295 83.495 104.465 ;
        RECT 83.785 104.295 83.955 104.465 ;
        RECT 84.245 104.295 84.415 104.465 ;
        RECT 84.705 104.295 84.875 104.465 ;
        RECT 85.165 104.295 85.335 104.465 ;
        RECT 85.625 104.295 85.795 104.465 ;
        RECT 86.085 104.295 86.255 104.465 ;
        RECT 86.545 104.295 86.715 104.465 ;
        RECT 87.005 104.295 87.175 104.465 ;
        RECT 87.465 104.295 87.635 104.465 ;
        RECT 87.925 104.295 88.095 104.465 ;
        RECT 88.385 104.295 88.555 104.465 ;
        RECT 88.845 104.295 89.015 104.465 ;
        RECT 89.305 104.295 89.475 104.465 ;
        RECT 89.765 104.295 89.935 104.465 ;
        RECT 90.225 104.295 90.395 104.465 ;
        RECT 90.685 104.295 90.855 104.465 ;
        RECT 91.145 104.295 91.315 104.465 ;
        RECT 91.605 104.295 91.775 104.465 ;
        RECT 92.065 104.295 92.235 104.465 ;
        RECT 92.525 104.295 92.695 104.465 ;
        RECT 92.985 104.295 93.155 104.465 ;
        RECT 93.445 104.295 93.615 104.465 ;
        RECT 93.905 104.295 94.075 104.465 ;
        RECT 94.365 104.295 94.535 104.465 ;
        RECT 94.825 104.295 94.995 104.465 ;
        RECT 95.285 104.295 95.455 104.465 ;
        RECT 95.745 104.295 95.915 104.465 ;
        RECT 96.205 104.295 96.375 104.465 ;
        RECT 96.665 104.295 96.835 104.465 ;
        RECT 97.125 104.295 97.295 104.465 ;
        RECT 97.585 104.295 97.755 104.465 ;
        RECT 98.045 104.295 98.215 104.465 ;
        RECT 98.505 104.295 98.675 104.465 ;
        RECT 98.965 104.295 99.135 104.465 ;
        RECT 99.425 104.295 99.595 104.465 ;
        RECT 99.885 104.295 100.055 104.465 ;
        RECT 100.345 104.295 100.515 104.465 ;
        RECT 100.805 104.295 100.975 104.465 ;
        RECT 101.265 104.295 101.435 104.465 ;
        RECT 101.725 104.295 101.895 104.465 ;
        RECT 102.185 104.295 102.355 104.465 ;
        RECT 102.645 104.295 102.815 104.465 ;
        RECT 103.105 104.295 103.275 104.465 ;
        RECT 103.565 104.295 103.735 104.465 ;
        RECT 104.025 104.295 104.195 104.465 ;
        RECT 104.485 104.295 104.655 104.465 ;
        RECT 104.945 104.295 105.115 104.465 ;
        RECT 105.405 104.295 105.575 104.465 ;
        RECT 105.865 104.295 106.035 104.465 ;
        RECT 106.325 104.295 106.495 104.465 ;
        RECT 106.785 104.295 106.955 104.465 ;
        RECT 107.245 104.295 107.415 104.465 ;
        RECT 107.705 104.295 107.875 104.465 ;
        RECT 108.165 104.295 108.335 104.465 ;
        RECT 108.625 104.295 108.795 104.465 ;
        RECT 109.085 104.295 109.255 104.465 ;
        RECT 109.545 104.295 109.715 104.465 ;
        RECT 110.005 104.295 110.175 104.465 ;
        RECT 110.465 104.295 110.635 104.465 ;
        RECT 110.925 104.295 111.095 104.465 ;
        RECT 111.385 104.295 111.555 104.465 ;
        RECT 111.845 104.295 112.015 104.465 ;
        RECT 112.305 104.295 112.475 104.465 ;
        RECT 112.765 104.295 112.935 104.465 ;
        RECT 113.225 104.295 113.395 104.465 ;
        RECT 113.685 104.295 113.855 104.465 ;
        RECT 114.145 104.295 114.315 104.465 ;
        RECT 114.605 104.295 114.775 104.465 ;
        RECT 115.065 104.295 115.235 104.465 ;
        RECT 115.525 104.295 115.695 104.465 ;
        RECT 115.985 104.295 116.155 104.465 ;
        RECT 116.445 104.295 116.615 104.465 ;
        RECT 116.905 104.295 117.075 104.465 ;
        RECT 117.365 104.295 117.535 104.465 ;
        RECT 117.825 104.295 117.995 104.465 ;
        RECT 118.285 104.295 118.455 104.465 ;
        RECT 118.745 104.295 118.915 104.465 ;
        RECT 119.205 104.295 119.375 104.465 ;
        RECT 119.665 104.295 119.835 104.465 ;
        RECT 120.125 104.295 120.295 104.465 ;
        RECT 120.585 104.295 120.755 104.465 ;
        RECT 121.045 104.295 121.215 104.465 ;
        RECT 121.505 104.295 121.675 104.465 ;
        RECT 121.965 104.295 122.135 104.465 ;
        RECT 122.425 104.295 122.595 104.465 ;
        RECT 122.885 104.295 123.055 104.465 ;
        RECT 123.345 104.295 123.515 104.465 ;
        RECT 123.805 104.295 123.975 104.465 ;
        RECT 124.265 104.295 124.435 104.465 ;
        RECT 124.725 104.295 124.895 104.465 ;
        RECT 125.185 104.295 125.355 104.465 ;
        RECT 125.645 104.295 125.815 104.465 ;
        RECT 126.105 104.295 126.275 104.465 ;
        RECT 126.565 104.295 126.735 104.465 ;
        RECT 127.025 104.295 127.195 104.465 ;
        RECT 127.485 104.295 127.655 104.465 ;
        RECT 127.945 104.295 128.115 104.465 ;
        RECT 128.405 104.295 128.575 104.465 ;
        RECT 128.865 104.295 129.035 104.465 ;
        RECT 129.325 104.295 129.495 104.465 ;
        RECT 129.785 104.295 129.955 104.465 ;
        RECT 130.245 104.295 130.415 104.465 ;
        RECT 130.705 104.295 130.875 104.465 ;
        RECT 131.165 104.295 131.335 104.465 ;
        RECT 131.625 104.295 131.795 104.465 ;
        RECT 132.085 104.295 132.255 104.465 ;
        RECT 132.545 104.295 132.715 104.465 ;
        RECT 133.005 104.295 133.175 104.465 ;
        RECT 133.465 104.295 133.635 104.465 ;
        RECT 133.925 104.295 134.095 104.465 ;
        RECT 134.385 104.295 134.555 104.465 ;
        RECT 134.845 104.295 135.015 104.465 ;
        RECT 135.305 104.295 135.475 104.465 ;
        RECT 135.765 104.295 135.935 104.465 ;
        RECT 136.225 104.295 136.395 104.465 ;
        RECT 136.685 104.295 136.855 104.465 ;
        RECT 137.145 104.295 137.315 104.465 ;
        RECT 137.605 104.295 137.775 104.465 ;
        RECT 138.065 104.295 138.235 104.465 ;
        RECT 138.525 104.295 138.695 104.465 ;
        RECT 138.985 104.295 139.155 104.465 ;
        RECT 52.965 103.785 53.135 103.955 ;
        RECT 52.045 103.105 52.215 103.275 ;
        RECT 61.705 103.445 61.875 103.615 ;
        RECT 59.865 103.105 60.035 103.275 ;
        RECT 61.245 103.105 61.415 103.275 ;
        RECT 62.170 103.105 62.340 103.275 ;
        RECT 63.085 103.445 63.255 103.615 ;
        RECT 65.400 103.105 65.570 103.275 ;
        RECT 62.625 102.765 62.795 102.935 ;
        RECT 64.005 102.765 64.175 102.935 ;
        RECT 50.665 101.575 50.835 101.745 ;
        RECT 51.125 101.575 51.295 101.745 ;
        RECT 51.585 101.575 51.755 101.745 ;
        RECT 52.045 101.575 52.215 101.745 ;
        RECT 52.505 101.575 52.675 101.745 ;
        RECT 52.965 101.575 53.135 101.745 ;
        RECT 53.425 101.575 53.595 101.745 ;
        RECT 53.885 101.575 54.055 101.745 ;
        RECT 54.345 101.575 54.515 101.745 ;
        RECT 54.805 101.575 54.975 101.745 ;
        RECT 55.265 101.575 55.435 101.745 ;
        RECT 55.725 101.575 55.895 101.745 ;
        RECT 56.185 101.575 56.355 101.745 ;
        RECT 56.645 101.575 56.815 101.745 ;
        RECT 57.105 101.575 57.275 101.745 ;
        RECT 57.565 101.575 57.735 101.745 ;
        RECT 58.025 101.575 58.195 101.745 ;
        RECT 58.485 101.575 58.655 101.745 ;
        RECT 58.945 101.575 59.115 101.745 ;
        RECT 59.405 101.575 59.575 101.745 ;
        RECT 59.865 101.575 60.035 101.745 ;
        RECT 60.325 101.575 60.495 101.745 ;
        RECT 60.785 101.575 60.955 101.745 ;
        RECT 61.245 101.575 61.415 101.745 ;
        RECT 61.705 101.575 61.875 101.745 ;
        RECT 62.165 101.575 62.335 101.745 ;
        RECT 62.625 101.575 62.795 101.745 ;
        RECT 63.085 101.575 63.255 101.745 ;
        RECT 63.545 101.575 63.715 101.745 ;
        RECT 64.005 101.575 64.175 101.745 ;
        RECT 64.465 101.575 64.635 101.745 ;
        RECT 64.925 101.575 65.095 101.745 ;
        RECT 65.385 101.575 65.555 101.745 ;
        RECT 65.845 101.575 66.015 101.745 ;
        RECT 66.305 101.575 66.475 101.745 ;
        RECT 66.765 101.575 66.935 101.745 ;
        RECT 67.225 101.575 67.395 101.745 ;
        RECT 67.685 101.575 67.855 101.745 ;
        RECT 68.145 101.575 68.315 101.745 ;
        RECT 68.605 101.575 68.775 101.745 ;
        RECT 69.065 101.575 69.235 101.745 ;
        RECT 69.525 101.575 69.695 101.745 ;
        RECT 69.985 101.575 70.155 101.745 ;
        RECT 70.445 101.575 70.615 101.745 ;
        RECT 70.905 101.575 71.075 101.745 ;
        RECT 71.365 101.575 71.535 101.745 ;
        RECT 71.825 101.575 71.995 101.745 ;
        RECT 72.285 101.575 72.455 101.745 ;
        RECT 72.745 101.575 72.915 101.745 ;
        RECT 73.205 101.575 73.375 101.745 ;
        RECT 73.665 101.575 73.835 101.745 ;
        RECT 74.125 101.575 74.295 101.745 ;
        RECT 74.585 101.575 74.755 101.745 ;
        RECT 75.045 101.575 75.215 101.745 ;
        RECT 75.505 101.575 75.675 101.745 ;
        RECT 75.965 101.575 76.135 101.745 ;
        RECT 76.425 101.575 76.595 101.745 ;
        RECT 76.885 101.575 77.055 101.745 ;
        RECT 77.345 101.575 77.515 101.745 ;
        RECT 77.805 101.575 77.975 101.745 ;
        RECT 78.265 101.575 78.435 101.745 ;
        RECT 78.725 101.575 78.895 101.745 ;
        RECT 79.185 101.575 79.355 101.745 ;
        RECT 79.645 101.575 79.815 101.745 ;
        RECT 80.105 101.575 80.275 101.745 ;
        RECT 80.565 101.575 80.735 101.745 ;
        RECT 81.025 101.575 81.195 101.745 ;
        RECT 81.485 101.575 81.655 101.745 ;
        RECT 81.945 101.575 82.115 101.745 ;
        RECT 82.405 101.575 82.575 101.745 ;
        RECT 82.865 101.575 83.035 101.745 ;
        RECT 83.325 101.575 83.495 101.745 ;
        RECT 83.785 101.575 83.955 101.745 ;
        RECT 84.245 101.575 84.415 101.745 ;
        RECT 84.705 101.575 84.875 101.745 ;
        RECT 85.165 101.575 85.335 101.745 ;
        RECT 85.625 101.575 85.795 101.745 ;
        RECT 86.085 101.575 86.255 101.745 ;
        RECT 86.545 101.575 86.715 101.745 ;
        RECT 87.005 101.575 87.175 101.745 ;
        RECT 87.465 101.575 87.635 101.745 ;
        RECT 87.925 101.575 88.095 101.745 ;
        RECT 88.385 101.575 88.555 101.745 ;
        RECT 88.845 101.575 89.015 101.745 ;
        RECT 89.305 101.575 89.475 101.745 ;
        RECT 89.765 101.575 89.935 101.745 ;
        RECT 90.225 101.575 90.395 101.745 ;
        RECT 90.685 101.575 90.855 101.745 ;
        RECT 91.145 101.575 91.315 101.745 ;
        RECT 91.605 101.575 91.775 101.745 ;
        RECT 92.065 101.575 92.235 101.745 ;
        RECT 92.525 101.575 92.695 101.745 ;
        RECT 92.985 101.575 93.155 101.745 ;
        RECT 93.445 101.575 93.615 101.745 ;
        RECT 93.905 101.575 94.075 101.745 ;
        RECT 94.365 101.575 94.535 101.745 ;
        RECT 94.825 101.575 94.995 101.745 ;
        RECT 95.285 101.575 95.455 101.745 ;
        RECT 95.745 101.575 95.915 101.745 ;
        RECT 96.205 101.575 96.375 101.745 ;
        RECT 96.665 101.575 96.835 101.745 ;
        RECT 97.125 101.575 97.295 101.745 ;
        RECT 97.585 101.575 97.755 101.745 ;
        RECT 98.045 101.575 98.215 101.745 ;
        RECT 98.505 101.575 98.675 101.745 ;
        RECT 98.965 101.575 99.135 101.745 ;
        RECT 99.425 101.575 99.595 101.745 ;
        RECT 99.885 101.575 100.055 101.745 ;
        RECT 100.345 101.575 100.515 101.745 ;
        RECT 100.805 101.575 100.975 101.745 ;
        RECT 101.265 101.575 101.435 101.745 ;
        RECT 101.725 101.575 101.895 101.745 ;
        RECT 102.185 101.575 102.355 101.745 ;
        RECT 102.645 101.575 102.815 101.745 ;
        RECT 103.105 101.575 103.275 101.745 ;
        RECT 103.565 101.575 103.735 101.745 ;
        RECT 104.025 101.575 104.195 101.745 ;
        RECT 104.485 101.575 104.655 101.745 ;
        RECT 104.945 101.575 105.115 101.745 ;
        RECT 105.405 101.575 105.575 101.745 ;
        RECT 105.865 101.575 106.035 101.745 ;
        RECT 106.325 101.575 106.495 101.745 ;
        RECT 106.785 101.575 106.955 101.745 ;
        RECT 107.245 101.575 107.415 101.745 ;
        RECT 107.705 101.575 107.875 101.745 ;
        RECT 108.165 101.575 108.335 101.745 ;
        RECT 108.625 101.575 108.795 101.745 ;
        RECT 109.085 101.575 109.255 101.745 ;
        RECT 109.545 101.575 109.715 101.745 ;
        RECT 110.005 101.575 110.175 101.745 ;
        RECT 110.465 101.575 110.635 101.745 ;
        RECT 110.925 101.575 111.095 101.745 ;
        RECT 111.385 101.575 111.555 101.745 ;
        RECT 111.845 101.575 112.015 101.745 ;
        RECT 112.305 101.575 112.475 101.745 ;
        RECT 112.765 101.575 112.935 101.745 ;
        RECT 113.225 101.575 113.395 101.745 ;
        RECT 113.685 101.575 113.855 101.745 ;
        RECT 114.145 101.575 114.315 101.745 ;
        RECT 114.605 101.575 114.775 101.745 ;
        RECT 115.065 101.575 115.235 101.745 ;
        RECT 115.525 101.575 115.695 101.745 ;
        RECT 115.985 101.575 116.155 101.745 ;
        RECT 116.445 101.575 116.615 101.745 ;
        RECT 116.905 101.575 117.075 101.745 ;
        RECT 117.365 101.575 117.535 101.745 ;
        RECT 117.825 101.575 117.995 101.745 ;
        RECT 118.285 101.575 118.455 101.745 ;
        RECT 118.745 101.575 118.915 101.745 ;
        RECT 119.205 101.575 119.375 101.745 ;
        RECT 119.665 101.575 119.835 101.745 ;
        RECT 120.125 101.575 120.295 101.745 ;
        RECT 120.585 101.575 120.755 101.745 ;
        RECT 121.045 101.575 121.215 101.745 ;
        RECT 121.505 101.575 121.675 101.745 ;
        RECT 121.965 101.575 122.135 101.745 ;
        RECT 122.425 101.575 122.595 101.745 ;
        RECT 122.885 101.575 123.055 101.745 ;
        RECT 123.345 101.575 123.515 101.745 ;
        RECT 123.805 101.575 123.975 101.745 ;
        RECT 124.265 101.575 124.435 101.745 ;
        RECT 124.725 101.575 124.895 101.745 ;
        RECT 125.185 101.575 125.355 101.745 ;
        RECT 125.645 101.575 125.815 101.745 ;
        RECT 126.105 101.575 126.275 101.745 ;
        RECT 126.565 101.575 126.735 101.745 ;
        RECT 127.025 101.575 127.195 101.745 ;
        RECT 127.485 101.575 127.655 101.745 ;
        RECT 127.945 101.575 128.115 101.745 ;
        RECT 128.405 101.575 128.575 101.745 ;
        RECT 128.865 101.575 129.035 101.745 ;
        RECT 129.325 101.575 129.495 101.745 ;
        RECT 129.785 101.575 129.955 101.745 ;
        RECT 130.245 101.575 130.415 101.745 ;
        RECT 130.705 101.575 130.875 101.745 ;
        RECT 131.165 101.575 131.335 101.745 ;
        RECT 131.625 101.575 131.795 101.745 ;
        RECT 132.085 101.575 132.255 101.745 ;
        RECT 132.545 101.575 132.715 101.745 ;
        RECT 133.005 101.575 133.175 101.745 ;
        RECT 133.465 101.575 133.635 101.745 ;
        RECT 133.925 101.575 134.095 101.745 ;
        RECT 134.385 101.575 134.555 101.745 ;
        RECT 134.845 101.575 135.015 101.745 ;
        RECT 135.305 101.575 135.475 101.745 ;
        RECT 135.765 101.575 135.935 101.745 ;
        RECT 136.225 101.575 136.395 101.745 ;
        RECT 136.685 101.575 136.855 101.745 ;
        RECT 137.145 101.575 137.315 101.745 ;
        RECT 137.605 101.575 137.775 101.745 ;
        RECT 138.065 101.575 138.235 101.745 ;
        RECT 138.525 101.575 138.695 101.745 ;
        RECT 138.985 101.575 139.155 101.745 ;
        RECT 52.045 100.045 52.215 100.215 ;
        RECT 52.965 99.365 53.135 99.535 ;
        RECT 50.665 98.855 50.835 99.025 ;
        RECT 51.125 98.855 51.295 99.025 ;
        RECT 51.585 98.855 51.755 99.025 ;
        RECT 52.045 98.855 52.215 99.025 ;
        RECT 52.505 98.855 52.675 99.025 ;
        RECT 52.965 98.855 53.135 99.025 ;
        RECT 53.425 98.855 53.595 99.025 ;
        RECT 53.885 98.855 54.055 99.025 ;
        RECT 54.345 98.855 54.515 99.025 ;
        RECT 54.805 98.855 54.975 99.025 ;
        RECT 55.265 98.855 55.435 99.025 ;
        RECT 55.725 98.855 55.895 99.025 ;
        RECT 56.185 98.855 56.355 99.025 ;
        RECT 56.645 98.855 56.815 99.025 ;
        RECT 57.105 98.855 57.275 99.025 ;
        RECT 57.565 98.855 57.735 99.025 ;
        RECT 58.025 98.855 58.195 99.025 ;
        RECT 58.485 98.855 58.655 99.025 ;
        RECT 58.945 98.855 59.115 99.025 ;
        RECT 59.405 98.855 59.575 99.025 ;
        RECT 59.865 98.855 60.035 99.025 ;
        RECT 60.325 98.855 60.495 99.025 ;
        RECT 60.785 98.855 60.955 99.025 ;
        RECT 61.245 98.855 61.415 99.025 ;
        RECT 61.705 98.855 61.875 99.025 ;
        RECT 62.165 98.855 62.335 99.025 ;
        RECT 62.625 98.855 62.795 99.025 ;
        RECT 63.085 98.855 63.255 99.025 ;
        RECT 63.545 98.855 63.715 99.025 ;
        RECT 64.005 98.855 64.175 99.025 ;
        RECT 64.465 98.855 64.635 99.025 ;
        RECT 64.925 98.855 65.095 99.025 ;
        RECT 65.385 98.855 65.555 99.025 ;
        RECT 65.845 98.855 66.015 99.025 ;
        RECT 66.305 98.855 66.475 99.025 ;
        RECT 66.765 98.855 66.935 99.025 ;
        RECT 67.225 98.855 67.395 99.025 ;
        RECT 67.685 98.855 67.855 99.025 ;
        RECT 68.145 98.855 68.315 99.025 ;
        RECT 68.605 98.855 68.775 99.025 ;
        RECT 69.065 98.855 69.235 99.025 ;
        RECT 69.525 98.855 69.695 99.025 ;
        RECT 69.985 98.855 70.155 99.025 ;
        RECT 70.445 98.855 70.615 99.025 ;
        RECT 70.905 98.855 71.075 99.025 ;
        RECT 71.365 98.855 71.535 99.025 ;
        RECT 71.825 98.855 71.995 99.025 ;
        RECT 72.285 98.855 72.455 99.025 ;
        RECT 72.745 98.855 72.915 99.025 ;
        RECT 73.205 98.855 73.375 99.025 ;
        RECT 73.665 98.855 73.835 99.025 ;
        RECT 74.125 98.855 74.295 99.025 ;
        RECT 74.585 98.855 74.755 99.025 ;
        RECT 75.045 98.855 75.215 99.025 ;
        RECT 75.505 98.855 75.675 99.025 ;
        RECT 75.965 98.855 76.135 99.025 ;
        RECT 76.425 98.855 76.595 99.025 ;
        RECT 76.885 98.855 77.055 99.025 ;
        RECT 77.345 98.855 77.515 99.025 ;
        RECT 77.805 98.855 77.975 99.025 ;
        RECT 78.265 98.855 78.435 99.025 ;
        RECT 78.725 98.855 78.895 99.025 ;
        RECT 79.185 98.855 79.355 99.025 ;
        RECT 79.645 98.855 79.815 99.025 ;
        RECT 80.105 98.855 80.275 99.025 ;
        RECT 80.565 98.855 80.735 99.025 ;
        RECT 81.025 98.855 81.195 99.025 ;
        RECT 81.485 98.855 81.655 99.025 ;
        RECT 81.945 98.855 82.115 99.025 ;
        RECT 82.405 98.855 82.575 99.025 ;
        RECT 82.865 98.855 83.035 99.025 ;
        RECT 83.325 98.855 83.495 99.025 ;
        RECT 83.785 98.855 83.955 99.025 ;
        RECT 84.245 98.855 84.415 99.025 ;
        RECT 84.705 98.855 84.875 99.025 ;
        RECT 85.165 98.855 85.335 99.025 ;
        RECT 85.625 98.855 85.795 99.025 ;
        RECT 86.085 98.855 86.255 99.025 ;
        RECT 86.545 98.855 86.715 99.025 ;
        RECT 87.005 98.855 87.175 99.025 ;
        RECT 87.465 98.855 87.635 99.025 ;
        RECT 87.925 98.855 88.095 99.025 ;
        RECT 88.385 98.855 88.555 99.025 ;
        RECT 88.845 98.855 89.015 99.025 ;
        RECT 89.305 98.855 89.475 99.025 ;
        RECT 89.765 98.855 89.935 99.025 ;
        RECT 90.225 98.855 90.395 99.025 ;
        RECT 90.685 98.855 90.855 99.025 ;
        RECT 91.145 98.855 91.315 99.025 ;
        RECT 91.605 98.855 91.775 99.025 ;
        RECT 92.065 98.855 92.235 99.025 ;
        RECT 92.525 98.855 92.695 99.025 ;
        RECT 92.985 98.855 93.155 99.025 ;
        RECT 93.445 98.855 93.615 99.025 ;
        RECT 93.905 98.855 94.075 99.025 ;
        RECT 94.365 98.855 94.535 99.025 ;
        RECT 94.825 98.855 94.995 99.025 ;
        RECT 95.285 98.855 95.455 99.025 ;
        RECT 95.745 98.855 95.915 99.025 ;
        RECT 96.205 98.855 96.375 99.025 ;
        RECT 96.665 98.855 96.835 99.025 ;
        RECT 97.125 98.855 97.295 99.025 ;
        RECT 97.585 98.855 97.755 99.025 ;
        RECT 98.045 98.855 98.215 99.025 ;
        RECT 98.505 98.855 98.675 99.025 ;
        RECT 98.965 98.855 99.135 99.025 ;
        RECT 99.425 98.855 99.595 99.025 ;
        RECT 99.885 98.855 100.055 99.025 ;
        RECT 100.345 98.855 100.515 99.025 ;
        RECT 100.805 98.855 100.975 99.025 ;
        RECT 101.265 98.855 101.435 99.025 ;
        RECT 101.725 98.855 101.895 99.025 ;
        RECT 102.185 98.855 102.355 99.025 ;
        RECT 102.645 98.855 102.815 99.025 ;
        RECT 103.105 98.855 103.275 99.025 ;
        RECT 103.565 98.855 103.735 99.025 ;
        RECT 104.025 98.855 104.195 99.025 ;
        RECT 104.485 98.855 104.655 99.025 ;
        RECT 104.945 98.855 105.115 99.025 ;
        RECT 105.405 98.855 105.575 99.025 ;
        RECT 105.865 98.855 106.035 99.025 ;
        RECT 106.325 98.855 106.495 99.025 ;
        RECT 106.785 98.855 106.955 99.025 ;
        RECT 107.245 98.855 107.415 99.025 ;
        RECT 107.705 98.855 107.875 99.025 ;
        RECT 108.165 98.855 108.335 99.025 ;
        RECT 108.625 98.855 108.795 99.025 ;
        RECT 109.085 98.855 109.255 99.025 ;
        RECT 109.545 98.855 109.715 99.025 ;
        RECT 110.005 98.855 110.175 99.025 ;
        RECT 110.465 98.855 110.635 99.025 ;
        RECT 110.925 98.855 111.095 99.025 ;
        RECT 111.385 98.855 111.555 99.025 ;
        RECT 111.845 98.855 112.015 99.025 ;
        RECT 112.305 98.855 112.475 99.025 ;
        RECT 112.765 98.855 112.935 99.025 ;
        RECT 113.225 98.855 113.395 99.025 ;
        RECT 113.685 98.855 113.855 99.025 ;
        RECT 114.145 98.855 114.315 99.025 ;
        RECT 114.605 98.855 114.775 99.025 ;
        RECT 115.065 98.855 115.235 99.025 ;
        RECT 115.525 98.855 115.695 99.025 ;
        RECT 115.985 98.855 116.155 99.025 ;
        RECT 116.445 98.855 116.615 99.025 ;
        RECT 116.905 98.855 117.075 99.025 ;
        RECT 117.365 98.855 117.535 99.025 ;
        RECT 117.825 98.855 117.995 99.025 ;
        RECT 118.285 98.855 118.455 99.025 ;
        RECT 118.745 98.855 118.915 99.025 ;
        RECT 119.205 98.855 119.375 99.025 ;
        RECT 119.665 98.855 119.835 99.025 ;
        RECT 120.125 98.855 120.295 99.025 ;
        RECT 120.585 98.855 120.755 99.025 ;
        RECT 121.045 98.855 121.215 99.025 ;
        RECT 121.505 98.855 121.675 99.025 ;
        RECT 121.965 98.855 122.135 99.025 ;
        RECT 122.425 98.855 122.595 99.025 ;
        RECT 122.885 98.855 123.055 99.025 ;
        RECT 123.345 98.855 123.515 99.025 ;
        RECT 123.805 98.855 123.975 99.025 ;
        RECT 124.265 98.855 124.435 99.025 ;
        RECT 124.725 98.855 124.895 99.025 ;
        RECT 125.185 98.855 125.355 99.025 ;
        RECT 125.645 98.855 125.815 99.025 ;
        RECT 126.105 98.855 126.275 99.025 ;
        RECT 126.565 98.855 126.735 99.025 ;
        RECT 127.025 98.855 127.195 99.025 ;
        RECT 127.485 98.855 127.655 99.025 ;
        RECT 127.945 98.855 128.115 99.025 ;
        RECT 128.405 98.855 128.575 99.025 ;
        RECT 128.865 98.855 129.035 99.025 ;
        RECT 129.325 98.855 129.495 99.025 ;
        RECT 129.785 98.855 129.955 99.025 ;
        RECT 130.245 98.855 130.415 99.025 ;
        RECT 130.705 98.855 130.875 99.025 ;
        RECT 131.165 98.855 131.335 99.025 ;
        RECT 131.625 98.855 131.795 99.025 ;
        RECT 132.085 98.855 132.255 99.025 ;
        RECT 132.545 98.855 132.715 99.025 ;
        RECT 133.005 98.855 133.175 99.025 ;
        RECT 133.465 98.855 133.635 99.025 ;
        RECT 133.925 98.855 134.095 99.025 ;
        RECT 134.385 98.855 134.555 99.025 ;
        RECT 134.845 98.855 135.015 99.025 ;
        RECT 135.305 98.855 135.475 99.025 ;
        RECT 135.765 98.855 135.935 99.025 ;
        RECT 136.225 98.855 136.395 99.025 ;
        RECT 136.685 98.855 136.855 99.025 ;
        RECT 137.145 98.855 137.315 99.025 ;
        RECT 137.605 98.855 137.775 99.025 ;
        RECT 138.065 98.855 138.235 99.025 ;
        RECT 138.525 98.855 138.695 99.025 ;
        RECT 138.985 98.855 139.155 99.025 ;
        RECT 61.705 98.345 61.875 98.515 ;
        RECT 60.785 97.665 60.955 97.835 ;
        RECT 50.665 96.135 50.835 96.305 ;
        RECT 51.125 96.135 51.295 96.305 ;
        RECT 51.585 96.135 51.755 96.305 ;
        RECT 52.045 96.135 52.215 96.305 ;
        RECT 52.505 96.135 52.675 96.305 ;
        RECT 52.965 96.135 53.135 96.305 ;
        RECT 53.425 96.135 53.595 96.305 ;
        RECT 53.885 96.135 54.055 96.305 ;
        RECT 54.345 96.135 54.515 96.305 ;
        RECT 54.805 96.135 54.975 96.305 ;
        RECT 55.265 96.135 55.435 96.305 ;
        RECT 55.725 96.135 55.895 96.305 ;
        RECT 56.185 96.135 56.355 96.305 ;
        RECT 56.645 96.135 56.815 96.305 ;
        RECT 57.105 96.135 57.275 96.305 ;
        RECT 57.565 96.135 57.735 96.305 ;
        RECT 58.025 96.135 58.195 96.305 ;
        RECT 58.485 96.135 58.655 96.305 ;
        RECT 58.945 96.135 59.115 96.305 ;
        RECT 59.405 96.135 59.575 96.305 ;
        RECT 59.865 96.135 60.035 96.305 ;
        RECT 60.325 96.135 60.495 96.305 ;
        RECT 60.785 96.135 60.955 96.305 ;
        RECT 61.245 96.135 61.415 96.305 ;
        RECT 61.705 96.135 61.875 96.305 ;
        RECT 62.165 96.135 62.335 96.305 ;
        RECT 62.625 96.135 62.795 96.305 ;
        RECT 63.085 96.135 63.255 96.305 ;
        RECT 63.545 96.135 63.715 96.305 ;
        RECT 64.005 96.135 64.175 96.305 ;
        RECT 64.465 96.135 64.635 96.305 ;
        RECT 64.925 96.135 65.095 96.305 ;
        RECT 65.385 96.135 65.555 96.305 ;
        RECT 65.845 96.135 66.015 96.305 ;
        RECT 66.305 96.135 66.475 96.305 ;
        RECT 66.765 96.135 66.935 96.305 ;
        RECT 67.225 96.135 67.395 96.305 ;
        RECT 67.685 96.135 67.855 96.305 ;
        RECT 68.145 96.135 68.315 96.305 ;
        RECT 68.605 96.135 68.775 96.305 ;
        RECT 69.065 96.135 69.235 96.305 ;
        RECT 69.525 96.135 69.695 96.305 ;
        RECT 69.985 96.135 70.155 96.305 ;
        RECT 70.445 96.135 70.615 96.305 ;
        RECT 70.905 96.135 71.075 96.305 ;
        RECT 71.365 96.135 71.535 96.305 ;
        RECT 71.825 96.135 71.995 96.305 ;
        RECT 72.285 96.135 72.455 96.305 ;
        RECT 72.745 96.135 72.915 96.305 ;
        RECT 73.205 96.135 73.375 96.305 ;
        RECT 73.665 96.135 73.835 96.305 ;
        RECT 74.125 96.135 74.295 96.305 ;
        RECT 74.585 96.135 74.755 96.305 ;
        RECT 75.045 96.135 75.215 96.305 ;
        RECT 75.505 96.135 75.675 96.305 ;
        RECT 75.965 96.135 76.135 96.305 ;
        RECT 76.425 96.135 76.595 96.305 ;
        RECT 76.885 96.135 77.055 96.305 ;
        RECT 77.345 96.135 77.515 96.305 ;
        RECT 77.805 96.135 77.975 96.305 ;
        RECT 78.265 96.135 78.435 96.305 ;
        RECT 78.725 96.135 78.895 96.305 ;
        RECT 79.185 96.135 79.355 96.305 ;
        RECT 79.645 96.135 79.815 96.305 ;
        RECT 80.105 96.135 80.275 96.305 ;
        RECT 80.565 96.135 80.735 96.305 ;
        RECT 81.025 96.135 81.195 96.305 ;
        RECT 81.485 96.135 81.655 96.305 ;
        RECT 81.945 96.135 82.115 96.305 ;
        RECT 82.405 96.135 82.575 96.305 ;
        RECT 82.865 96.135 83.035 96.305 ;
        RECT 83.325 96.135 83.495 96.305 ;
        RECT 83.785 96.135 83.955 96.305 ;
        RECT 84.245 96.135 84.415 96.305 ;
        RECT 84.705 96.135 84.875 96.305 ;
        RECT 85.165 96.135 85.335 96.305 ;
        RECT 85.625 96.135 85.795 96.305 ;
        RECT 86.085 96.135 86.255 96.305 ;
        RECT 86.545 96.135 86.715 96.305 ;
        RECT 87.005 96.135 87.175 96.305 ;
        RECT 87.465 96.135 87.635 96.305 ;
        RECT 87.925 96.135 88.095 96.305 ;
        RECT 88.385 96.135 88.555 96.305 ;
        RECT 88.845 96.135 89.015 96.305 ;
        RECT 89.305 96.135 89.475 96.305 ;
        RECT 89.765 96.135 89.935 96.305 ;
        RECT 90.225 96.135 90.395 96.305 ;
        RECT 90.685 96.135 90.855 96.305 ;
        RECT 91.145 96.135 91.315 96.305 ;
        RECT 91.605 96.135 91.775 96.305 ;
        RECT 92.065 96.135 92.235 96.305 ;
        RECT 92.525 96.135 92.695 96.305 ;
        RECT 92.985 96.135 93.155 96.305 ;
        RECT 93.445 96.135 93.615 96.305 ;
        RECT 93.905 96.135 94.075 96.305 ;
        RECT 94.365 96.135 94.535 96.305 ;
        RECT 94.825 96.135 94.995 96.305 ;
        RECT 95.285 96.135 95.455 96.305 ;
        RECT 95.745 96.135 95.915 96.305 ;
        RECT 96.205 96.135 96.375 96.305 ;
        RECT 96.665 96.135 96.835 96.305 ;
        RECT 97.125 96.135 97.295 96.305 ;
        RECT 97.585 96.135 97.755 96.305 ;
        RECT 98.045 96.135 98.215 96.305 ;
        RECT 98.505 96.135 98.675 96.305 ;
        RECT 98.965 96.135 99.135 96.305 ;
        RECT 99.425 96.135 99.595 96.305 ;
        RECT 99.885 96.135 100.055 96.305 ;
        RECT 100.345 96.135 100.515 96.305 ;
        RECT 100.805 96.135 100.975 96.305 ;
        RECT 101.265 96.135 101.435 96.305 ;
        RECT 101.725 96.135 101.895 96.305 ;
        RECT 102.185 96.135 102.355 96.305 ;
        RECT 102.645 96.135 102.815 96.305 ;
        RECT 103.105 96.135 103.275 96.305 ;
        RECT 103.565 96.135 103.735 96.305 ;
        RECT 104.025 96.135 104.195 96.305 ;
        RECT 104.485 96.135 104.655 96.305 ;
        RECT 104.945 96.135 105.115 96.305 ;
        RECT 105.405 96.135 105.575 96.305 ;
        RECT 105.865 96.135 106.035 96.305 ;
        RECT 106.325 96.135 106.495 96.305 ;
        RECT 106.785 96.135 106.955 96.305 ;
        RECT 107.245 96.135 107.415 96.305 ;
        RECT 107.705 96.135 107.875 96.305 ;
        RECT 108.165 96.135 108.335 96.305 ;
        RECT 108.625 96.135 108.795 96.305 ;
        RECT 109.085 96.135 109.255 96.305 ;
        RECT 109.545 96.135 109.715 96.305 ;
        RECT 110.005 96.135 110.175 96.305 ;
        RECT 110.465 96.135 110.635 96.305 ;
        RECT 110.925 96.135 111.095 96.305 ;
        RECT 111.385 96.135 111.555 96.305 ;
        RECT 111.845 96.135 112.015 96.305 ;
        RECT 112.305 96.135 112.475 96.305 ;
        RECT 112.765 96.135 112.935 96.305 ;
        RECT 113.225 96.135 113.395 96.305 ;
        RECT 113.685 96.135 113.855 96.305 ;
        RECT 114.145 96.135 114.315 96.305 ;
        RECT 114.605 96.135 114.775 96.305 ;
        RECT 115.065 96.135 115.235 96.305 ;
        RECT 115.525 96.135 115.695 96.305 ;
        RECT 115.985 96.135 116.155 96.305 ;
        RECT 116.445 96.135 116.615 96.305 ;
        RECT 116.905 96.135 117.075 96.305 ;
        RECT 117.365 96.135 117.535 96.305 ;
        RECT 117.825 96.135 117.995 96.305 ;
        RECT 118.285 96.135 118.455 96.305 ;
        RECT 118.745 96.135 118.915 96.305 ;
        RECT 119.205 96.135 119.375 96.305 ;
        RECT 119.665 96.135 119.835 96.305 ;
        RECT 120.125 96.135 120.295 96.305 ;
        RECT 120.585 96.135 120.755 96.305 ;
        RECT 121.045 96.135 121.215 96.305 ;
        RECT 121.505 96.135 121.675 96.305 ;
        RECT 121.965 96.135 122.135 96.305 ;
        RECT 122.425 96.135 122.595 96.305 ;
        RECT 122.885 96.135 123.055 96.305 ;
        RECT 123.345 96.135 123.515 96.305 ;
        RECT 123.805 96.135 123.975 96.305 ;
        RECT 124.265 96.135 124.435 96.305 ;
        RECT 124.725 96.135 124.895 96.305 ;
        RECT 125.185 96.135 125.355 96.305 ;
        RECT 125.645 96.135 125.815 96.305 ;
        RECT 126.105 96.135 126.275 96.305 ;
        RECT 126.565 96.135 126.735 96.305 ;
        RECT 127.025 96.135 127.195 96.305 ;
        RECT 127.485 96.135 127.655 96.305 ;
        RECT 127.945 96.135 128.115 96.305 ;
        RECT 128.405 96.135 128.575 96.305 ;
        RECT 128.865 96.135 129.035 96.305 ;
        RECT 129.325 96.135 129.495 96.305 ;
        RECT 129.785 96.135 129.955 96.305 ;
        RECT 130.245 96.135 130.415 96.305 ;
        RECT 130.705 96.135 130.875 96.305 ;
        RECT 131.165 96.135 131.335 96.305 ;
        RECT 131.625 96.135 131.795 96.305 ;
        RECT 132.085 96.135 132.255 96.305 ;
        RECT 132.545 96.135 132.715 96.305 ;
        RECT 133.005 96.135 133.175 96.305 ;
        RECT 133.465 96.135 133.635 96.305 ;
        RECT 133.925 96.135 134.095 96.305 ;
        RECT 134.385 96.135 134.555 96.305 ;
        RECT 134.845 96.135 135.015 96.305 ;
        RECT 135.305 96.135 135.475 96.305 ;
        RECT 135.765 96.135 135.935 96.305 ;
        RECT 136.225 96.135 136.395 96.305 ;
        RECT 136.685 96.135 136.855 96.305 ;
        RECT 137.145 96.135 137.315 96.305 ;
        RECT 137.605 96.135 137.775 96.305 ;
        RECT 138.065 96.135 138.235 96.305 ;
        RECT 138.525 96.135 138.695 96.305 ;
        RECT 138.985 96.135 139.155 96.305 ;
        RECT 61.705 94.605 61.875 94.775 ;
        RECT 62.625 94.605 62.795 94.775 ;
        RECT 61.705 93.925 61.875 94.095 ;
        RECT 50.665 93.415 50.835 93.585 ;
        RECT 51.125 93.415 51.295 93.585 ;
        RECT 51.585 93.415 51.755 93.585 ;
        RECT 52.045 93.415 52.215 93.585 ;
        RECT 52.505 93.415 52.675 93.585 ;
        RECT 52.965 93.415 53.135 93.585 ;
        RECT 53.425 93.415 53.595 93.585 ;
        RECT 53.885 93.415 54.055 93.585 ;
        RECT 54.345 93.415 54.515 93.585 ;
        RECT 54.805 93.415 54.975 93.585 ;
        RECT 55.265 93.415 55.435 93.585 ;
        RECT 55.725 93.415 55.895 93.585 ;
        RECT 56.185 93.415 56.355 93.585 ;
        RECT 56.645 93.415 56.815 93.585 ;
        RECT 57.105 93.415 57.275 93.585 ;
        RECT 57.565 93.415 57.735 93.585 ;
        RECT 58.025 93.415 58.195 93.585 ;
        RECT 58.485 93.415 58.655 93.585 ;
        RECT 58.945 93.415 59.115 93.585 ;
        RECT 59.405 93.415 59.575 93.585 ;
        RECT 59.865 93.415 60.035 93.585 ;
        RECT 60.325 93.415 60.495 93.585 ;
        RECT 60.785 93.415 60.955 93.585 ;
        RECT 61.245 93.415 61.415 93.585 ;
        RECT 61.705 93.415 61.875 93.585 ;
        RECT 62.165 93.415 62.335 93.585 ;
        RECT 62.625 93.415 62.795 93.585 ;
        RECT 63.085 93.415 63.255 93.585 ;
        RECT 63.545 93.415 63.715 93.585 ;
        RECT 64.005 93.415 64.175 93.585 ;
        RECT 64.465 93.415 64.635 93.585 ;
        RECT 64.925 93.415 65.095 93.585 ;
        RECT 65.385 93.415 65.555 93.585 ;
        RECT 65.845 93.415 66.015 93.585 ;
        RECT 66.305 93.415 66.475 93.585 ;
        RECT 66.765 93.415 66.935 93.585 ;
        RECT 67.225 93.415 67.395 93.585 ;
        RECT 67.685 93.415 67.855 93.585 ;
        RECT 68.145 93.415 68.315 93.585 ;
        RECT 68.605 93.415 68.775 93.585 ;
        RECT 69.065 93.415 69.235 93.585 ;
        RECT 69.525 93.415 69.695 93.585 ;
        RECT 69.985 93.415 70.155 93.585 ;
        RECT 70.445 93.415 70.615 93.585 ;
        RECT 70.905 93.415 71.075 93.585 ;
        RECT 71.365 93.415 71.535 93.585 ;
        RECT 71.825 93.415 71.995 93.585 ;
        RECT 72.285 93.415 72.455 93.585 ;
        RECT 72.745 93.415 72.915 93.585 ;
        RECT 73.205 93.415 73.375 93.585 ;
        RECT 73.665 93.415 73.835 93.585 ;
        RECT 74.125 93.415 74.295 93.585 ;
        RECT 74.585 93.415 74.755 93.585 ;
        RECT 75.045 93.415 75.215 93.585 ;
        RECT 75.505 93.415 75.675 93.585 ;
        RECT 75.965 93.415 76.135 93.585 ;
        RECT 76.425 93.415 76.595 93.585 ;
        RECT 76.885 93.415 77.055 93.585 ;
        RECT 77.345 93.415 77.515 93.585 ;
        RECT 77.805 93.415 77.975 93.585 ;
        RECT 78.265 93.415 78.435 93.585 ;
        RECT 78.725 93.415 78.895 93.585 ;
        RECT 79.185 93.415 79.355 93.585 ;
        RECT 79.645 93.415 79.815 93.585 ;
        RECT 80.105 93.415 80.275 93.585 ;
        RECT 80.565 93.415 80.735 93.585 ;
        RECT 81.025 93.415 81.195 93.585 ;
        RECT 81.485 93.415 81.655 93.585 ;
        RECT 81.945 93.415 82.115 93.585 ;
        RECT 82.405 93.415 82.575 93.585 ;
        RECT 82.865 93.415 83.035 93.585 ;
        RECT 83.325 93.415 83.495 93.585 ;
        RECT 83.785 93.415 83.955 93.585 ;
        RECT 84.245 93.415 84.415 93.585 ;
        RECT 84.705 93.415 84.875 93.585 ;
        RECT 85.165 93.415 85.335 93.585 ;
        RECT 85.625 93.415 85.795 93.585 ;
        RECT 86.085 93.415 86.255 93.585 ;
        RECT 86.545 93.415 86.715 93.585 ;
        RECT 87.005 93.415 87.175 93.585 ;
        RECT 87.465 93.415 87.635 93.585 ;
        RECT 87.925 93.415 88.095 93.585 ;
        RECT 88.385 93.415 88.555 93.585 ;
        RECT 88.845 93.415 89.015 93.585 ;
        RECT 89.305 93.415 89.475 93.585 ;
        RECT 89.765 93.415 89.935 93.585 ;
        RECT 90.225 93.415 90.395 93.585 ;
        RECT 90.685 93.415 90.855 93.585 ;
        RECT 91.145 93.415 91.315 93.585 ;
        RECT 91.605 93.415 91.775 93.585 ;
        RECT 92.065 93.415 92.235 93.585 ;
        RECT 92.525 93.415 92.695 93.585 ;
        RECT 92.985 93.415 93.155 93.585 ;
        RECT 93.445 93.415 93.615 93.585 ;
        RECT 93.905 93.415 94.075 93.585 ;
        RECT 94.365 93.415 94.535 93.585 ;
        RECT 94.825 93.415 94.995 93.585 ;
        RECT 95.285 93.415 95.455 93.585 ;
        RECT 95.745 93.415 95.915 93.585 ;
        RECT 96.205 93.415 96.375 93.585 ;
        RECT 96.665 93.415 96.835 93.585 ;
        RECT 97.125 93.415 97.295 93.585 ;
        RECT 97.585 93.415 97.755 93.585 ;
        RECT 98.045 93.415 98.215 93.585 ;
        RECT 98.505 93.415 98.675 93.585 ;
        RECT 98.965 93.415 99.135 93.585 ;
        RECT 99.425 93.415 99.595 93.585 ;
        RECT 99.885 93.415 100.055 93.585 ;
        RECT 100.345 93.415 100.515 93.585 ;
        RECT 100.805 93.415 100.975 93.585 ;
        RECT 101.265 93.415 101.435 93.585 ;
        RECT 101.725 93.415 101.895 93.585 ;
        RECT 102.185 93.415 102.355 93.585 ;
        RECT 102.645 93.415 102.815 93.585 ;
        RECT 103.105 93.415 103.275 93.585 ;
        RECT 103.565 93.415 103.735 93.585 ;
        RECT 104.025 93.415 104.195 93.585 ;
        RECT 104.485 93.415 104.655 93.585 ;
        RECT 104.945 93.415 105.115 93.585 ;
        RECT 105.405 93.415 105.575 93.585 ;
        RECT 105.865 93.415 106.035 93.585 ;
        RECT 106.325 93.415 106.495 93.585 ;
        RECT 106.785 93.415 106.955 93.585 ;
        RECT 107.245 93.415 107.415 93.585 ;
        RECT 107.705 93.415 107.875 93.585 ;
        RECT 108.165 93.415 108.335 93.585 ;
        RECT 108.625 93.415 108.795 93.585 ;
        RECT 109.085 93.415 109.255 93.585 ;
        RECT 109.545 93.415 109.715 93.585 ;
        RECT 110.005 93.415 110.175 93.585 ;
        RECT 110.465 93.415 110.635 93.585 ;
        RECT 110.925 93.415 111.095 93.585 ;
        RECT 111.385 93.415 111.555 93.585 ;
        RECT 111.845 93.415 112.015 93.585 ;
        RECT 112.305 93.415 112.475 93.585 ;
        RECT 112.765 93.415 112.935 93.585 ;
        RECT 113.225 93.415 113.395 93.585 ;
        RECT 113.685 93.415 113.855 93.585 ;
        RECT 114.145 93.415 114.315 93.585 ;
        RECT 114.605 93.415 114.775 93.585 ;
        RECT 115.065 93.415 115.235 93.585 ;
        RECT 115.525 93.415 115.695 93.585 ;
        RECT 115.985 93.415 116.155 93.585 ;
        RECT 116.445 93.415 116.615 93.585 ;
        RECT 116.905 93.415 117.075 93.585 ;
        RECT 117.365 93.415 117.535 93.585 ;
        RECT 117.825 93.415 117.995 93.585 ;
        RECT 118.285 93.415 118.455 93.585 ;
        RECT 118.745 93.415 118.915 93.585 ;
        RECT 119.205 93.415 119.375 93.585 ;
        RECT 119.665 93.415 119.835 93.585 ;
        RECT 120.125 93.415 120.295 93.585 ;
        RECT 120.585 93.415 120.755 93.585 ;
        RECT 121.045 93.415 121.215 93.585 ;
        RECT 121.505 93.415 121.675 93.585 ;
        RECT 121.965 93.415 122.135 93.585 ;
        RECT 122.425 93.415 122.595 93.585 ;
        RECT 122.885 93.415 123.055 93.585 ;
        RECT 123.345 93.415 123.515 93.585 ;
        RECT 123.805 93.415 123.975 93.585 ;
        RECT 124.265 93.415 124.435 93.585 ;
        RECT 124.725 93.415 124.895 93.585 ;
        RECT 125.185 93.415 125.355 93.585 ;
        RECT 125.645 93.415 125.815 93.585 ;
        RECT 126.105 93.415 126.275 93.585 ;
        RECT 126.565 93.415 126.735 93.585 ;
        RECT 127.025 93.415 127.195 93.585 ;
        RECT 127.485 93.415 127.655 93.585 ;
        RECT 127.945 93.415 128.115 93.585 ;
        RECT 128.405 93.415 128.575 93.585 ;
        RECT 128.865 93.415 129.035 93.585 ;
        RECT 129.325 93.415 129.495 93.585 ;
        RECT 129.785 93.415 129.955 93.585 ;
        RECT 130.245 93.415 130.415 93.585 ;
        RECT 130.705 93.415 130.875 93.585 ;
        RECT 131.165 93.415 131.335 93.585 ;
        RECT 131.625 93.415 131.795 93.585 ;
        RECT 132.085 93.415 132.255 93.585 ;
        RECT 132.545 93.415 132.715 93.585 ;
        RECT 133.005 93.415 133.175 93.585 ;
        RECT 133.465 93.415 133.635 93.585 ;
        RECT 133.925 93.415 134.095 93.585 ;
        RECT 134.385 93.415 134.555 93.585 ;
        RECT 134.845 93.415 135.015 93.585 ;
        RECT 135.305 93.415 135.475 93.585 ;
        RECT 135.765 93.415 135.935 93.585 ;
        RECT 136.225 93.415 136.395 93.585 ;
        RECT 136.685 93.415 136.855 93.585 ;
        RECT 137.145 93.415 137.315 93.585 ;
        RECT 137.605 93.415 137.775 93.585 ;
        RECT 138.065 93.415 138.235 93.585 ;
        RECT 138.525 93.415 138.695 93.585 ;
        RECT 138.985 93.415 139.155 93.585 ;
        RECT 58.025 92.905 58.195 93.075 ;
        RECT 57.565 91.885 57.735 92.055 ;
        RECT 58.485 92.905 58.655 93.075 ;
        RECT 60.325 91.205 60.495 91.375 ;
        RECT 60.785 92.905 60.955 93.075 ;
        RECT 63.085 92.565 63.255 92.735 ;
        RECT 63.545 91.885 63.715 92.055 ;
        RECT 64.925 92.225 65.095 92.395 ;
        RECT 66.765 92.565 66.935 92.735 ;
        RECT 66.305 92.225 66.475 92.395 ;
        RECT 50.665 90.695 50.835 90.865 ;
        RECT 51.125 90.695 51.295 90.865 ;
        RECT 51.585 90.695 51.755 90.865 ;
        RECT 52.045 90.695 52.215 90.865 ;
        RECT 52.505 90.695 52.675 90.865 ;
        RECT 52.965 90.695 53.135 90.865 ;
        RECT 53.425 90.695 53.595 90.865 ;
        RECT 53.885 90.695 54.055 90.865 ;
        RECT 54.345 90.695 54.515 90.865 ;
        RECT 54.805 90.695 54.975 90.865 ;
        RECT 55.265 90.695 55.435 90.865 ;
        RECT 55.725 90.695 55.895 90.865 ;
        RECT 56.185 90.695 56.355 90.865 ;
        RECT 56.645 90.695 56.815 90.865 ;
        RECT 57.105 90.695 57.275 90.865 ;
        RECT 57.565 90.695 57.735 90.865 ;
        RECT 58.025 90.695 58.195 90.865 ;
        RECT 58.485 90.695 58.655 90.865 ;
        RECT 58.945 90.695 59.115 90.865 ;
        RECT 59.405 90.695 59.575 90.865 ;
        RECT 59.865 90.695 60.035 90.865 ;
        RECT 60.325 90.695 60.495 90.865 ;
        RECT 60.785 90.695 60.955 90.865 ;
        RECT 61.245 90.695 61.415 90.865 ;
        RECT 61.705 90.695 61.875 90.865 ;
        RECT 62.165 90.695 62.335 90.865 ;
        RECT 62.625 90.695 62.795 90.865 ;
        RECT 63.085 90.695 63.255 90.865 ;
        RECT 63.545 90.695 63.715 90.865 ;
        RECT 64.005 90.695 64.175 90.865 ;
        RECT 64.465 90.695 64.635 90.865 ;
        RECT 64.925 90.695 65.095 90.865 ;
        RECT 65.385 90.695 65.555 90.865 ;
        RECT 65.845 90.695 66.015 90.865 ;
        RECT 66.305 90.695 66.475 90.865 ;
        RECT 66.765 90.695 66.935 90.865 ;
        RECT 67.225 90.695 67.395 90.865 ;
        RECT 67.685 90.695 67.855 90.865 ;
        RECT 68.145 90.695 68.315 90.865 ;
        RECT 68.605 90.695 68.775 90.865 ;
        RECT 69.065 90.695 69.235 90.865 ;
        RECT 69.525 90.695 69.695 90.865 ;
        RECT 69.985 90.695 70.155 90.865 ;
        RECT 70.445 90.695 70.615 90.865 ;
        RECT 70.905 90.695 71.075 90.865 ;
        RECT 71.365 90.695 71.535 90.865 ;
        RECT 71.825 90.695 71.995 90.865 ;
        RECT 72.285 90.695 72.455 90.865 ;
        RECT 72.745 90.695 72.915 90.865 ;
        RECT 73.205 90.695 73.375 90.865 ;
        RECT 73.665 90.695 73.835 90.865 ;
        RECT 74.125 90.695 74.295 90.865 ;
        RECT 74.585 90.695 74.755 90.865 ;
        RECT 75.045 90.695 75.215 90.865 ;
        RECT 75.505 90.695 75.675 90.865 ;
        RECT 75.965 90.695 76.135 90.865 ;
        RECT 76.425 90.695 76.595 90.865 ;
        RECT 76.885 90.695 77.055 90.865 ;
        RECT 77.345 90.695 77.515 90.865 ;
        RECT 77.805 90.695 77.975 90.865 ;
        RECT 78.265 90.695 78.435 90.865 ;
        RECT 78.725 90.695 78.895 90.865 ;
        RECT 79.185 90.695 79.355 90.865 ;
        RECT 79.645 90.695 79.815 90.865 ;
        RECT 80.105 90.695 80.275 90.865 ;
        RECT 80.565 90.695 80.735 90.865 ;
        RECT 81.025 90.695 81.195 90.865 ;
        RECT 81.485 90.695 81.655 90.865 ;
        RECT 81.945 90.695 82.115 90.865 ;
        RECT 82.405 90.695 82.575 90.865 ;
        RECT 82.865 90.695 83.035 90.865 ;
        RECT 83.325 90.695 83.495 90.865 ;
        RECT 83.785 90.695 83.955 90.865 ;
        RECT 84.245 90.695 84.415 90.865 ;
        RECT 84.705 90.695 84.875 90.865 ;
        RECT 85.165 90.695 85.335 90.865 ;
        RECT 85.625 90.695 85.795 90.865 ;
        RECT 86.085 90.695 86.255 90.865 ;
        RECT 86.545 90.695 86.715 90.865 ;
        RECT 87.005 90.695 87.175 90.865 ;
        RECT 87.465 90.695 87.635 90.865 ;
        RECT 87.925 90.695 88.095 90.865 ;
        RECT 88.385 90.695 88.555 90.865 ;
        RECT 88.845 90.695 89.015 90.865 ;
        RECT 89.305 90.695 89.475 90.865 ;
        RECT 89.765 90.695 89.935 90.865 ;
        RECT 90.225 90.695 90.395 90.865 ;
        RECT 90.685 90.695 90.855 90.865 ;
        RECT 91.145 90.695 91.315 90.865 ;
        RECT 91.605 90.695 91.775 90.865 ;
        RECT 92.065 90.695 92.235 90.865 ;
        RECT 92.525 90.695 92.695 90.865 ;
        RECT 92.985 90.695 93.155 90.865 ;
        RECT 93.445 90.695 93.615 90.865 ;
        RECT 93.905 90.695 94.075 90.865 ;
        RECT 94.365 90.695 94.535 90.865 ;
        RECT 94.825 90.695 94.995 90.865 ;
        RECT 95.285 90.695 95.455 90.865 ;
        RECT 95.745 90.695 95.915 90.865 ;
        RECT 96.205 90.695 96.375 90.865 ;
        RECT 96.665 90.695 96.835 90.865 ;
        RECT 97.125 90.695 97.295 90.865 ;
        RECT 97.585 90.695 97.755 90.865 ;
        RECT 98.045 90.695 98.215 90.865 ;
        RECT 98.505 90.695 98.675 90.865 ;
        RECT 98.965 90.695 99.135 90.865 ;
        RECT 99.425 90.695 99.595 90.865 ;
        RECT 99.885 90.695 100.055 90.865 ;
        RECT 100.345 90.695 100.515 90.865 ;
        RECT 100.805 90.695 100.975 90.865 ;
        RECT 101.265 90.695 101.435 90.865 ;
        RECT 101.725 90.695 101.895 90.865 ;
        RECT 102.185 90.695 102.355 90.865 ;
        RECT 102.645 90.695 102.815 90.865 ;
        RECT 103.105 90.695 103.275 90.865 ;
        RECT 103.565 90.695 103.735 90.865 ;
        RECT 104.025 90.695 104.195 90.865 ;
        RECT 104.485 90.695 104.655 90.865 ;
        RECT 104.945 90.695 105.115 90.865 ;
        RECT 105.405 90.695 105.575 90.865 ;
        RECT 105.865 90.695 106.035 90.865 ;
        RECT 106.325 90.695 106.495 90.865 ;
        RECT 106.785 90.695 106.955 90.865 ;
        RECT 107.245 90.695 107.415 90.865 ;
        RECT 107.705 90.695 107.875 90.865 ;
        RECT 108.165 90.695 108.335 90.865 ;
        RECT 108.625 90.695 108.795 90.865 ;
        RECT 109.085 90.695 109.255 90.865 ;
        RECT 109.545 90.695 109.715 90.865 ;
        RECT 110.005 90.695 110.175 90.865 ;
        RECT 110.465 90.695 110.635 90.865 ;
        RECT 110.925 90.695 111.095 90.865 ;
        RECT 111.385 90.695 111.555 90.865 ;
        RECT 111.845 90.695 112.015 90.865 ;
        RECT 112.305 90.695 112.475 90.865 ;
        RECT 112.765 90.695 112.935 90.865 ;
        RECT 113.225 90.695 113.395 90.865 ;
        RECT 113.685 90.695 113.855 90.865 ;
        RECT 114.145 90.695 114.315 90.865 ;
        RECT 114.605 90.695 114.775 90.865 ;
        RECT 115.065 90.695 115.235 90.865 ;
        RECT 115.525 90.695 115.695 90.865 ;
        RECT 115.985 90.695 116.155 90.865 ;
        RECT 116.445 90.695 116.615 90.865 ;
        RECT 116.905 90.695 117.075 90.865 ;
        RECT 117.365 90.695 117.535 90.865 ;
        RECT 117.825 90.695 117.995 90.865 ;
        RECT 118.285 90.695 118.455 90.865 ;
        RECT 118.745 90.695 118.915 90.865 ;
        RECT 119.205 90.695 119.375 90.865 ;
        RECT 119.665 90.695 119.835 90.865 ;
        RECT 120.125 90.695 120.295 90.865 ;
        RECT 120.585 90.695 120.755 90.865 ;
        RECT 121.045 90.695 121.215 90.865 ;
        RECT 121.505 90.695 121.675 90.865 ;
        RECT 121.965 90.695 122.135 90.865 ;
        RECT 122.425 90.695 122.595 90.865 ;
        RECT 122.885 90.695 123.055 90.865 ;
        RECT 123.345 90.695 123.515 90.865 ;
        RECT 123.805 90.695 123.975 90.865 ;
        RECT 124.265 90.695 124.435 90.865 ;
        RECT 124.725 90.695 124.895 90.865 ;
        RECT 125.185 90.695 125.355 90.865 ;
        RECT 125.645 90.695 125.815 90.865 ;
        RECT 126.105 90.695 126.275 90.865 ;
        RECT 126.565 90.695 126.735 90.865 ;
        RECT 127.025 90.695 127.195 90.865 ;
        RECT 127.485 90.695 127.655 90.865 ;
        RECT 127.945 90.695 128.115 90.865 ;
        RECT 128.405 90.695 128.575 90.865 ;
        RECT 128.865 90.695 129.035 90.865 ;
        RECT 129.325 90.695 129.495 90.865 ;
        RECT 129.785 90.695 129.955 90.865 ;
        RECT 130.245 90.695 130.415 90.865 ;
        RECT 130.705 90.695 130.875 90.865 ;
        RECT 131.165 90.695 131.335 90.865 ;
        RECT 131.625 90.695 131.795 90.865 ;
        RECT 132.085 90.695 132.255 90.865 ;
        RECT 132.545 90.695 132.715 90.865 ;
        RECT 133.005 90.695 133.175 90.865 ;
        RECT 133.465 90.695 133.635 90.865 ;
        RECT 133.925 90.695 134.095 90.865 ;
        RECT 134.385 90.695 134.555 90.865 ;
        RECT 134.845 90.695 135.015 90.865 ;
        RECT 135.305 90.695 135.475 90.865 ;
        RECT 135.765 90.695 135.935 90.865 ;
        RECT 136.225 90.695 136.395 90.865 ;
        RECT 136.685 90.695 136.855 90.865 ;
        RECT 137.145 90.695 137.315 90.865 ;
        RECT 137.605 90.695 137.775 90.865 ;
        RECT 138.065 90.695 138.235 90.865 ;
        RECT 138.525 90.695 138.695 90.865 ;
        RECT 138.985 90.695 139.155 90.865 ;
        RECT 60.325 89.165 60.495 89.335 ;
        RECT 62.165 90.185 62.335 90.355 ;
        RECT 61.705 89.165 61.875 89.335 ;
        RECT 50.665 87.975 50.835 88.145 ;
        RECT 51.125 87.975 51.295 88.145 ;
        RECT 51.585 87.975 51.755 88.145 ;
        RECT 52.045 87.975 52.215 88.145 ;
        RECT 52.505 87.975 52.675 88.145 ;
        RECT 52.965 87.975 53.135 88.145 ;
        RECT 53.425 87.975 53.595 88.145 ;
        RECT 53.885 87.975 54.055 88.145 ;
        RECT 54.345 87.975 54.515 88.145 ;
        RECT 54.805 87.975 54.975 88.145 ;
        RECT 55.265 87.975 55.435 88.145 ;
        RECT 55.725 87.975 55.895 88.145 ;
        RECT 56.185 87.975 56.355 88.145 ;
        RECT 56.645 87.975 56.815 88.145 ;
        RECT 57.105 87.975 57.275 88.145 ;
        RECT 57.565 87.975 57.735 88.145 ;
        RECT 58.025 87.975 58.195 88.145 ;
        RECT 58.485 87.975 58.655 88.145 ;
        RECT 58.945 87.975 59.115 88.145 ;
        RECT 59.405 87.975 59.575 88.145 ;
        RECT 59.865 87.975 60.035 88.145 ;
        RECT 60.325 87.975 60.495 88.145 ;
        RECT 60.785 87.975 60.955 88.145 ;
        RECT 61.245 87.975 61.415 88.145 ;
        RECT 61.705 87.975 61.875 88.145 ;
        RECT 62.165 87.975 62.335 88.145 ;
        RECT 62.625 87.975 62.795 88.145 ;
        RECT 63.085 87.975 63.255 88.145 ;
        RECT 63.545 87.975 63.715 88.145 ;
        RECT 64.005 87.975 64.175 88.145 ;
        RECT 64.465 87.975 64.635 88.145 ;
        RECT 64.925 87.975 65.095 88.145 ;
        RECT 65.385 87.975 65.555 88.145 ;
        RECT 65.845 87.975 66.015 88.145 ;
        RECT 66.305 87.975 66.475 88.145 ;
        RECT 66.765 87.975 66.935 88.145 ;
        RECT 67.225 87.975 67.395 88.145 ;
        RECT 67.685 87.975 67.855 88.145 ;
        RECT 68.145 87.975 68.315 88.145 ;
        RECT 68.605 87.975 68.775 88.145 ;
        RECT 69.065 87.975 69.235 88.145 ;
        RECT 69.525 87.975 69.695 88.145 ;
        RECT 69.985 87.975 70.155 88.145 ;
        RECT 70.445 87.975 70.615 88.145 ;
        RECT 70.905 87.975 71.075 88.145 ;
        RECT 71.365 87.975 71.535 88.145 ;
        RECT 71.825 87.975 71.995 88.145 ;
        RECT 72.285 87.975 72.455 88.145 ;
        RECT 72.745 87.975 72.915 88.145 ;
        RECT 73.205 87.975 73.375 88.145 ;
        RECT 73.665 87.975 73.835 88.145 ;
        RECT 74.125 87.975 74.295 88.145 ;
        RECT 74.585 87.975 74.755 88.145 ;
        RECT 75.045 87.975 75.215 88.145 ;
        RECT 75.505 87.975 75.675 88.145 ;
        RECT 75.965 87.975 76.135 88.145 ;
        RECT 76.425 87.975 76.595 88.145 ;
        RECT 76.885 87.975 77.055 88.145 ;
        RECT 77.345 87.975 77.515 88.145 ;
        RECT 77.805 87.975 77.975 88.145 ;
        RECT 78.265 87.975 78.435 88.145 ;
        RECT 78.725 87.975 78.895 88.145 ;
        RECT 79.185 87.975 79.355 88.145 ;
        RECT 79.645 87.975 79.815 88.145 ;
        RECT 80.105 87.975 80.275 88.145 ;
        RECT 80.565 87.975 80.735 88.145 ;
        RECT 81.025 87.975 81.195 88.145 ;
        RECT 81.485 87.975 81.655 88.145 ;
        RECT 81.945 87.975 82.115 88.145 ;
        RECT 82.405 87.975 82.575 88.145 ;
        RECT 82.865 87.975 83.035 88.145 ;
        RECT 83.325 87.975 83.495 88.145 ;
        RECT 83.785 87.975 83.955 88.145 ;
        RECT 84.245 87.975 84.415 88.145 ;
        RECT 84.705 87.975 84.875 88.145 ;
        RECT 85.165 87.975 85.335 88.145 ;
        RECT 85.625 87.975 85.795 88.145 ;
        RECT 86.085 87.975 86.255 88.145 ;
        RECT 86.545 87.975 86.715 88.145 ;
        RECT 87.005 87.975 87.175 88.145 ;
        RECT 87.465 87.975 87.635 88.145 ;
        RECT 87.925 87.975 88.095 88.145 ;
        RECT 88.385 87.975 88.555 88.145 ;
        RECT 88.845 87.975 89.015 88.145 ;
        RECT 89.305 87.975 89.475 88.145 ;
        RECT 89.765 87.975 89.935 88.145 ;
        RECT 90.225 87.975 90.395 88.145 ;
        RECT 90.685 87.975 90.855 88.145 ;
        RECT 91.145 87.975 91.315 88.145 ;
        RECT 91.605 87.975 91.775 88.145 ;
        RECT 92.065 87.975 92.235 88.145 ;
        RECT 92.525 87.975 92.695 88.145 ;
        RECT 92.985 87.975 93.155 88.145 ;
        RECT 93.445 87.975 93.615 88.145 ;
        RECT 93.905 87.975 94.075 88.145 ;
        RECT 94.365 87.975 94.535 88.145 ;
        RECT 94.825 87.975 94.995 88.145 ;
        RECT 95.285 87.975 95.455 88.145 ;
        RECT 95.745 87.975 95.915 88.145 ;
        RECT 96.205 87.975 96.375 88.145 ;
        RECT 96.665 87.975 96.835 88.145 ;
        RECT 97.125 87.975 97.295 88.145 ;
        RECT 97.585 87.975 97.755 88.145 ;
        RECT 98.045 87.975 98.215 88.145 ;
        RECT 98.505 87.975 98.675 88.145 ;
        RECT 98.965 87.975 99.135 88.145 ;
        RECT 99.425 87.975 99.595 88.145 ;
        RECT 99.885 87.975 100.055 88.145 ;
        RECT 100.345 87.975 100.515 88.145 ;
        RECT 100.805 87.975 100.975 88.145 ;
        RECT 101.265 87.975 101.435 88.145 ;
        RECT 101.725 87.975 101.895 88.145 ;
        RECT 102.185 87.975 102.355 88.145 ;
        RECT 102.645 87.975 102.815 88.145 ;
        RECT 103.105 87.975 103.275 88.145 ;
        RECT 103.565 87.975 103.735 88.145 ;
        RECT 104.025 87.975 104.195 88.145 ;
        RECT 104.485 87.975 104.655 88.145 ;
        RECT 104.945 87.975 105.115 88.145 ;
        RECT 105.405 87.975 105.575 88.145 ;
        RECT 105.865 87.975 106.035 88.145 ;
        RECT 106.325 87.975 106.495 88.145 ;
        RECT 106.785 87.975 106.955 88.145 ;
        RECT 107.245 87.975 107.415 88.145 ;
        RECT 107.705 87.975 107.875 88.145 ;
        RECT 108.165 87.975 108.335 88.145 ;
        RECT 108.625 87.975 108.795 88.145 ;
        RECT 109.085 87.975 109.255 88.145 ;
        RECT 109.545 87.975 109.715 88.145 ;
        RECT 110.005 87.975 110.175 88.145 ;
        RECT 110.465 87.975 110.635 88.145 ;
        RECT 110.925 87.975 111.095 88.145 ;
        RECT 111.385 87.975 111.555 88.145 ;
        RECT 111.845 87.975 112.015 88.145 ;
        RECT 112.305 87.975 112.475 88.145 ;
        RECT 112.765 87.975 112.935 88.145 ;
        RECT 113.225 87.975 113.395 88.145 ;
        RECT 113.685 87.975 113.855 88.145 ;
        RECT 114.145 87.975 114.315 88.145 ;
        RECT 114.605 87.975 114.775 88.145 ;
        RECT 115.065 87.975 115.235 88.145 ;
        RECT 115.525 87.975 115.695 88.145 ;
        RECT 115.985 87.975 116.155 88.145 ;
        RECT 116.445 87.975 116.615 88.145 ;
        RECT 116.905 87.975 117.075 88.145 ;
        RECT 117.365 87.975 117.535 88.145 ;
        RECT 117.825 87.975 117.995 88.145 ;
        RECT 118.285 87.975 118.455 88.145 ;
        RECT 118.745 87.975 118.915 88.145 ;
        RECT 119.205 87.975 119.375 88.145 ;
        RECT 119.665 87.975 119.835 88.145 ;
        RECT 120.125 87.975 120.295 88.145 ;
        RECT 120.585 87.975 120.755 88.145 ;
        RECT 121.045 87.975 121.215 88.145 ;
        RECT 121.505 87.975 121.675 88.145 ;
        RECT 121.965 87.975 122.135 88.145 ;
        RECT 122.425 87.975 122.595 88.145 ;
        RECT 122.885 87.975 123.055 88.145 ;
        RECT 123.345 87.975 123.515 88.145 ;
        RECT 123.805 87.975 123.975 88.145 ;
        RECT 124.265 87.975 124.435 88.145 ;
        RECT 124.725 87.975 124.895 88.145 ;
        RECT 125.185 87.975 125.355 88.145 ;
        RECT 125.645 87.975 125.815 88.145 ;
        RECT 126.105 87.975 126.275 88.145 ;
        RECT 126.565 87.975 126.735 88.145 ;
        RECT 127.025 87.975 127.195 88.145 ;
        RECT 127.485 87.975 127.655 88.145 ;
        RECT 127.945 87.975 128.115 88.145 ;
        RECT 128.405 87.975 128.575 88.145 ;
        RECT 128.865 87.975 129.035 88.145 ;
        RECT 129.325 87.975 129.495 88.145 ;
        RECT 129.785 87.975 129.955 88.145 ;
        RECT 130.245 87.975 130.415 88.145 ;
        RECT 130.705 87.975 130.875 88.145 ;
        RECT 131.165 87.975 131.335 88.145 ;
        RECT 131.625 87.975 131.795 88.145 ;
        RECT 132.085 87.975 132.255 88.145 ;
        RECT 132.545 87.975 132.715 88.145 ;
        RECT 133.005 87.975 133.175 88.145 ;
        RECT 133.465 87.975 133.635 88.145 ;
        RECT 133.925 87.975 134.095 88.145 ;
        RECT 134.385 87.975 134.555 88.145 ;
        RECT 134.845 87.975 135.015 88.145 ;
        RECT 135.305 87.975 135.475 88.145 ;
        RECT 135.765 87.975 135.935 88.145 ;
        RECT 136.225 87.975 136.395 88.145 ;
        RECT 136.685 87.975 136.855 88.145 ;
        RECT 137.145 87.975 137.315 88.145 ;
        RECT 137.605 87.975 137.775 88.145 ;
        RECT 138.065 87.975 138.235 88.145 ;
        RECT 138.525 87.975 138.695 88.145 ;
        RECT 138.985 87.975 139.155 88.145 ;
        RECT 50.665 85.255 50.835 85.425 ;
        RECT 51.125 85.255 51.295 85.425 ;
        RECT 51.585 85.255 51.755 85.425 ;
        RECT 52.045 85.255 52.215 85.425 ;
        RECT 52.505 85.255 52.675 85.425 ;
        RECT 52.965 85.255 53.135 85.425 ;
        RECT 53.425 85.255 53.595 85.425 ;
        RECT 53.885 85.255 54.055 85.425 ;
        RECT 54.345 85.255 54.515 85.425 ;
        RECT 54.805 85.255 54.975 85.425 ;
        RECT 55.265 85.255 55.435 85.425 ;
        RECT 55.725 85.255 55.895 85.425 ;
        RECT 56.185 85.255 56.355 85.425 ;
        RECT 56.645 85.255 56.815 85.425 ;
        RECT 57.105 85.255 57.275 85.425 ;
        RECT 57.565 85.255 57.735 85.425 ;
        RECT 58.025 85.255 58.195 85.425 ;
        RECT 58.485 85.255 58.655 85.425 ;
        RECT 58.945 85.255 59.115 85.425 ;
        RECT 59.405 85.255 59.575 85.425 ;
        RECT 59.865 85.255 60.035 85.425 ;
        RECT 60.325 85.255 60.495 85.425 ;
        RECT 60.785 85.255 60.955 85.425 ;
        RECT 61.245 85.255 61.415 85.425 ;
        RECT 61.705 85.255 61.875 85.425 ;
        RECT 62.165 85.255 62.335 85.425 ;
        RECT 62.625 85.255 62.795 85.425 ;
        RECT 63.085 85.255 63.255 85.425 ;
        RECT 63.545 85.255 63.715 85.425 ;
        RECT 64.005 85.255 64.175 85.425 ;
        RECT 64.465 85.255 64.635 85.425 ;
        RECT 64.925 85.255 65.095 85.425 ;
        RECT 65.385 85.255 65.555 85.425 ;
        RECT 65.845 85.255 66.015 85.425 ;
        RECT 66.305 85.255 66.475 85.425 ;
        RECT 66.765 85.255 66.935 85.425 ;
        RECT 67.225 85.255 67.395 85.425 ;
        RECT 67.685 85.255 67.855 85.425 ;
        RECT 68.145 85.255 68.315 85.425 ;
        RECT 68.605 85.255 68.775 85.425 ;
        RECT 69.065 85.255 69.235 85.425 ;
        RECT 69.525 85.255 69.695 85.425 ;
        RECT 69.985 85.255 70.155 85.425 ;
        RECT 70.445 85.255 70.615 85.425 ;
        RECT 70.905 85.255 71.075 85.425 ;
        RECT 71.365 85.255 71.535 85.425 ;
        RECT 71.825 85.255 71.995 85.425 ;
        RECT 72.285 85.255 72.455 85.425 ;
        RECT 72.745 85.255 72.915 85.425 ;
        RECT 73.205 85.255 73.375 85.425 ;
        RECT 73.665 85.255 73.835 85.425 ;
        RECT 74.125 85.255 74.295 85.425 ;
        RECT 74.585 85.255 74.755 85.425 ;
        RECT 75.045 85.255 75.215 85.425 ;
        RECT 75.505 85.255 75.675 85.425 ;
        RECT 75.965 85.255 76.135 85.425 ;
        RECT 76.425 85.255 76.595 85.425 ;
        RECT 76.885 85.255 77.055 85.425 ;
        RECT 77.345 85.255 77.515 85.425 ;
        RECT 77.805 85.255 77.975 85.425 ;
        RECT 78.265 85.255 78.435 85.425 ;
        RECT 78.725 85.255 78.895 85.425 ;
        RECT 79.185 85.255 79.355 85.425 ;
        RECT 79.645 85.255 79.815 85.425 ;
        RECT 80.105 85.255 80.275 85.425 ;
        RECT 80.565 85.255 80.735 85.425 ;
        RECT 81.025 85.255 81.195 85.425 ;
        RECT 81.485 85.255 81.655 85.425 ;
        RECT 81.945 85.255 82.115 85.425 ;
        RECT 82.405 85.255 82.575 85.425 ;
        RECT 82.865 85.255 83.035 85.425 ;
        RECT 83.325 85.255 83.495 85.425 ;
        RECT 83.785 85.255 83.955 85.425 ;
        RECT 84.245 85.255 84.415 85.425 ;
        RECT 84.705 85.255 84.875 85.425 ;
        RECT 85.165 85.255 85.335 85.425 ;
        RECT 85.625 85.255 85.795 85.425 ;
        RECT 86.085 85.255 86.255 85.425 ;
        RECT 86.545 85.255 86.715 85.425 ;
        RECT 87.005 85.255 87.175 85.425 ;
        RECT 87.465 85.255 87.635 85.425 ;
        RECT 87.925 85.255 88.095 85.425 ;
        RECT 88.385 85.255 88.555 85.425 ;
        RECT 88.845 85.255 89.015 85.425 ;
        RECT 89.305 85.255 89.475 85.425 ;
        RECT 89.765 85.255 89.935 85.425 ;
        RECT 90.225 85.255 90.395 85.425 ;
        RECT 90.685 85.255 90.855 85.425 ;
        RECT 91.145 85.255 91.315 85.425 ;
        RECT 91.605 85.255 91.775 85.425 ;
        RECT 92.065 85.255 92.235 85.425 ;
        RECT 92.525 85.255 92.695 85.425 ;
        RECT 92.985 85.255 93.155 85.425 ;
        RECT 93.445 85.255 93.615 85.425 ;
        RECT 93.905 85.255 94.075 85.425 ;
        RECT 94.365 85.255 94.535 85.425 ;
        RECT 94.825 85.255 94.995 85.425 ;
        RECT 95.285 85.255 95.455 85.425 ;
        RECT 95.745 85.255 95.915 85.425 ;
        RECT 96.205 85.255 96.375 85.425 ;
        RECT 96.665 85.255 96.835 85.425 ;
        RECT 97.125 85.255 97.295 85.425 ;
        RECT 97.585 85.255 97.755 85.425 ;
        RECT 98.045 85.255 98.215 85.425 ;
        RECT 98.505 85.255 98.675 85.425 ;
        RECT 98.965 85.255 99.135 85.425 ;
        RECT 99.425 85.255 99.595 85.425 ;
        RECT 99.885 85.255 100.055 85.425 ;
        RECT 100.345 85.255 100.515 85.425 ;
        RECT 100.805 85.255 100.975 85.425 ;
        RECT 101.265 85.255 101.435 85.425 ;
        RECT 101.725 85.255 101.895 85.425 ;
        RECT 102.185 85.255 102.355 85.425 ;
        RECT 102.645 85.255 102.815 85.425 ;
        RECT 103.105 85.255 103.275 85.425 ;
        RECT 103.565 85.255 103.735 85.425 ;
        RECT 104.025 85.255 104.195 85.425 ;
        RECT 104.485 85.255 104.655 85.425 ;
        RECT 104.945 85.255 105.115 85.425 ;
        RECT 105.405 85.255 105.575 85.425 ;
        RECT 105.865 85.255 106.035 85.425 ;
        RECT 106.325 85.255 106.495 85.425 ;
        RECT 106.785 85.255 106.955 85.425 ;
        RECT 107.245 85.255 107.415 85.425 ;
        RECT 107.705 85.255 107.875 85.425 ;
        RECT 108.165 85.255 108.335 85.425 ;
        RECT 108.625 85.255 108.795 85.425 ;
        RECT 109.085 85.255 109.255 85.425 ;
        RECT 109.545 85.255 109.715 85.425 ;
        RECT 110.005 85.255 110.175 85.425 ;
        RECT 110.465 85.255 110.635 85.425 ;
        RECT 110.925 85.255 111.095 85.425 ;
        RECT 111.385 85.255 111.555 85.425 ;
        RECT 111.845 85.255 112.015 85.425 ;
        RECT 112.305 85.255 112.475 85.425 ;
        RECT 112.765 85.255 112.935 85.425 ;
        RECT 113.225 85.255 113.395 85.425 ;
        RECT 113.685 85.255 113.855 85.425 ;
        RECT 114.145 85.255 114.315 85.425 ;
        RECT 114.605 85.255 114.775 85.425 ;
        RECT 115.065 85.255 115.235 85.425 ;
        RECT 115.525 85.255 115.695 85.425 ;
        RECT 115.985 85.255 116.155 85.425 ;
        RECT 116.445 85.255 116.615 85.425 ;
        RECT 116.905 85.255 117.075 85.425 ;
        RECT 117.365 85.255 117.535 85.425 ;
        RECT 117.825 85.255 117.995 85.425 ;
        RECT 118.285 85.255 118.455 85.425 ;
        RECT 118.745 85.255 118.915 85.425 ;
        RECT 119.205 85.255 119.375 85.425 ;
        RECT 119.665 85.255 119.835 85.425 ;
        RECT 120.125 85.255 120.295 85.425 ;
        RECT 120.585 85.255 120.755 85.425 ;
        RECT 121.045 85.255 121.215 85.425 ;
        RECT 121.505 85.255 121.675 85.425 ;
        RECT 121.965 85.255 122.135 85.425 ;
        RECT 122.425 85.255 122.595 85.425 ;
        RECT 122.885 85.255 123.055 85.425 ;
        RECT 123.345 85.255 123.515 85.425 ;
        RECT 123.805 85.255 123.975 85.425 ;
        RECT 124.265 85.255 124.435 85.425 ;
        RECT 124.725 85.255 124.895 85.425 ;
        RECT 125.185 85.255 125.355 85.425 ;
        RECT 125.645 85.255 125.815 85.425 ;
        RECT 126.105 85.255 126.275 85.425 ;
        RECT 126.565 85.255 126.735 85.425 ;
        RECT 127.025 85.255 127.195 85.425 ;
        RECT 127.485 85.255 127.655 85.425 ;
        RECT 127.945 85.255 128.115 85.425 ;
        RECT 128.405 85.255 128.575 85.425 ;
        RECT 128.865 85.255 129.035 85.425 ;
        RECT 129.325 85.255 129.495 85.425 ;
        RECT 129.785 85.255 129.955 85.425 ;
        RECT 130.245 85.255 130.415 85.425 ;
        RECT 130.705 85.255 130.875 85.425 ;
        RECT 131.165 85.255 131.335 85.425 ;
        RECT 131.625 85.255 131.795 85.425 ;
        RECT 132.085 85.255 132.255 85.425 ;
        RECT 132.545 85.255 132.715 85.425 ;
        RECT 133.005 85.255 133.175 85.425 ;
        RECT 133.465 85.255 133.635 85.425 ;
        RECT 133.925 85.255 134.095 85.425 ;
        RECT 134.385 85.255 134.555 85.425 ;
        RECT 134.845 85.255 135.015 85.425 ;
        RECT 135.305 85.255 135.475 85.425 ;
        RECT 135.765 85.255 135.935 85.425 ;
        RECT 136.225 85.255 136.395 85.425 ;
        RECT 136.685 85.255 136.855 85.425 ;
        RECT 137.145 85.255 137.315 85.425 ;
        RECT 137.605 85.255 137.775 85.425 ;
        RECT 138.065 85.255 138.235 85.425 ;
        RECT 138.525 85.255 138.695 85.425 ;
        RECT 138.985 85.255 139.155 85.425 ;
        RECT 50.665 82.535 50.835 82.705 ;
        RECT 51.125 82.535 51.295 82.705 ;
        RECT 51.585 82.535 51.755 82.705 ;
        RECT 52.045 82.535 52.215 82.705 ;
        RECT 52.505 82.535 52.675 82.705 ;
        RECT 52.965 82.535 53.135 82.705 ;
        RECT 53.425 82.535 53.595 82.705 ;
        RECT 53.885 82.535 54.055 82.705 ;
        RECT 54.345 82.535 54.515 82.705 ;
        RECT 54.805 82.535 54.975 82.705 ;
        RECT 55.265 82.535 55.435 82.705 ;
        RECT 55.725 82.535 55.895 82.705 ;
        RECT 56.185 82.535 56.355 82.705 ;
        RECT 56.645 82.535 56.815 82.705 ;
        RECT 57.105 82.535 57.275 82.705 ;
        RECT 57.565 82.535 57.735 82.705 ;
        RECT 58.025 82.535 58.195 82.705 ;
        RECT 58.485 82.535 58.655 82.705 ;
        RECT 58.945 82.535 59.115 82.705 ;
        RECT 59.405 82.535 59.575 82.705 ;
        RECT 59.865 82.535 60.035 82.705 ;
        RECT 60.325 82.535 60.495 82.705 ;
        RECT 60.785 82.535 60.955 82.705 ;
        RECT 61.245 82.535 61.415 82.705 ;
        RECT 61.705 82.535 61.875 82.705 ;
        RECT 62.165 82.535 62.335 82.705 ;
        RECT 62.625 82.535 62.795 82.705 ;
        RECT 63.085 82.535 63.255 82.705 ;
        RECT 63.545 82.535 63.715 82.705 ;
        RECT 64.005 82.535 64.175 82.705 ;
        RECT 64.465 82.535 64.635 82.705 ;
        RECT 64.925 82.535 65.095 82.705 ;
        RECT 65.385 82.535 65.555 82.705 ;
        RECT 65.845 82.535 66.015 82.705 ;
        RECT 66.305 82.535 66.475 82.705 ;
        RECT 66.765 82.535 66.935 82.705 ;
        RECT 67.225 82.535 67.395 82.705 ;
        RECT 67.685 82.535 67.855 82.705 ;
        RECT 68.145 82.535 68.315 82.705 ;
        RECT 68.605 82.535 68.775 82.705 ;
        RECT 69.065 82.535 69.235 82.705 ;
        RECT 69.525 82.535 69.695 82.705 ;
        RECT 69.985 82.535 70.155 82.705 ;
        RECT 70.445 82.535 70.615 82.705 ;
        RECT 70.905 82.535 71.075 82.705 ;
        RECT 71.365 82.535 71.535 82.705 ;
        RECT 71.825 82.535 71.995 82.705 ;
        RECT 72.285 82.535 72.455 82.705 ;
        RECT 72.745 82.535 72.915 82.705 ;
        RECT 73.205 82.535 73.375 82.705 ;
        RECT 73.665 82.535 73.835 82.705 ;
        RECT 74.125 82.535 74.295 82.705 ;
        RECT 74.585 82.535 74.755 82.705 ;
        RECT 75.045 82.535 75.215 82.705 ;
        RECT 75.505 82.535 75.675 82.705 ;
        RECT 75.965 82.535 76.135 82.705 ;
        RECT 76.425 82.535 76.595 82.705 ;
        RECT 76.885 82.535 77.055 82.705 ;
        RECT 77.345 82.535 77.515 82.705 ;
        RECT 77.805 82.535 77.975 82.705 ;
        RECT 78.265 82.535 78.435 82.705 ;
        RECT 78.725 82.535 78.895 82.705 ;
        RECT 79.185 82.535 79.355 82.705 ;
        RECT 79.645 82.535 79.815 82.705 ;
        RECT 80.105 82.535 80.275 82.705 ;
        RECT 80.565 82.535 80.735 82.705 ;
        RECT 81.025 82.535 81.195 82.705 ;
        RECT 81.485 82.535 81.655 82.705 ;
        RECT 81.945 82.535 82.115 82.705 ;
        RECT 82.405 82.535 82.575 82.705 ;
        RECT 82.865 82.535 83.035 82.705 ;
        RECT 83.325 82.535 83.495 82.705 ;
        RECT 83.785 82.535 83.955 82.705 ;
        RECT 84.245 82.535 84.415 82.705 ;
        RECT 84.705 82.535 84.875 82.705 ;
        RECT 85.165 82.535 85.335 82.705 ;
        RECT 85.625 82.535 85.795 82.705 ;
        RECT 86.085 82.535 86.255 82.705 ;
        RECT 86.545 82.535 86.715 82.705 ;
        RECT 87.005 82.535 87.175 82.705 ;
        RECT 87.465 82.535 87.635 82.705 ;
        RECT 87.925 82.535 88.095 82.705 ;
        RECT 88.385 82.535 88.555 82.705 ;
        RECT 88.845 82.535 89.015 82.705 ;
        RECT 89.305 82.535 89.475 82.705 ;
        RECT 89.765 82.535 89.935 82.705 ;
        RECT 90.225 82.535 90.395 82.705 ;
        RECT 90.685 82.535 90.855 82.705 ;
        RECT 91.145 82.535 91.315 82.705 ;
        RECT 91.605 82.535 91.775 82.705 ;
        RECT 92.065 82.535 92.235 82.705 ;
        RECT 92.525 82.535 92.695 82.705 ;
        RECT 92.985 82.535 93.155 82.705 ;
        RECT 93.445 82.535 93.615 82.705 ;
        RECT 93.905 82.535 94.075 82.705 ;
        RECT 94.365 82.535 94.535 82.705 ;
        RECT 94.825 82.535 94.995 82.705 ;
        RECT 95.285 82.535 95.455 82.705 ;
        RECT 95.745 82.535 95.915 82.705 ;
        RECT 96.205 82.535 96.375 82.705 ;
        RECT 96.665 82.535 96.835 82.705 ;
        RECT 97.125 82.535 97.295 82.705 ;
        RECT 97.585 82.535 97.755 82.705 ;
        RECT 98.045 82.535 98.215 82.705 ;
        RECT 98.505 82.535 98.675 82.705 ;
        RECT 98.965 82.535 99.135 82.705 ;
        RECT 99.425 82.535 99.595 82.705 ;
        RECT 99.885 82.535 100.055 82.705 ;
        RECT 100.345 82.535 100.515 82.705 ;
        RECT 100.805 82.535 100.975 82.705 ;
        RECT 101.265 82.535 101.435 82.705 ;
        RECT 101.725 82.535 101.895 82.705 ;
        RECT 102.185 82.535 102.355 82.705 ;
        RECT 102.645 82.535 102.815 82.705 ;
        RECT 103.105 82.535 103.275 82.705 ;
        RECT 103.565 82.535 103.735 82.705 ;
        RECT 104.025 82.535 104.195 82.705 ;
        RECT 104.485 82.535 104.655 82.705 ;
        RECT 104.945 82.535 105.115 82.705 ;
        RECT 105.405 82.535 105.575 82.705 ;
        RECT 105.865 82.535 106.035 82.705 ;
        RECT 106.325 82.535 106.495 82.705 ;
        RECT 106.785 82.535 106.955 82.705 ;
        RECT 107.245 82.535 107.415 82.705 ;
        RECT 107.705 82.535 107.875 82.705 ;
        RECT 108.165 82.535 108.335 82.705 ;
        RECT 108.625 82.535 108.795 82.705 ;
        RECT 109.085 82.535 109.255 82.705 ;
        RECT 109.545 82.535 109.715 82.705 ;
        RECT 110.005 82.535 110.175 82.705 ;
        RECT 110.465 82.535 110.635 82.705 ;
        RECT 110.925 82.535 111.095 82.705 ;
        RECT 111.385 82.535 111.555 82.705 ;
        RECT 111.845 82.535 112.015 82.705 ;
        RECT 112.305 82.535 112.475 82.705 ;
        RECT 112.765 82.535 112.935 82.705 ;
        RECT 113.225 82.535 113.395 82.705 ;
        RECT 113.685 82.535 113.855 82.705 ;
        RECT 114.145 82.535 114.315 82.705 ;
        RECT 114.605 82.535 114.775 82.705 ;
        RECT 115.065 82.535 115.235 82.705 ;
        RECT 115.525 82.535 115.695 82.705 ;
        RECT 115.985 82.535 116.155 82.705 ;
        RECT 116.445 82.535 116.615 82.705 ;
        RECT 116.905 82.535 117.075 82.705 ;
        RECT 117.365 82.535 117.535 82.705 ;
        RECT 117.825 82.535 117.995 82.705 ;
        RECT 118.285 82.535 118.455 82.705 ;
        RECT 118.745 82.535 118.915 82.705 ;
        RECT 119.205 82.535 119.375 82.705 ;
        RECT 119.665 82.535 119.835 82.705 ;
        RECT 120.125 82.535 120.295 82.705 ;
        RECT 120.585 82.535 120.755 82.705 ;
        RECT 121.045 82.535 121.215 82.705 ;
        RECT 121.505 82.535 121.675 82.705 ;
        RECT 121.965 82.535 122.135 82.705 ;
        RECT 122.425 82.535 122.595 82.705 ;
        RECT 122.885 82.535 123.055 82.705 ;
        RECT 123.345 82.535 123.515 82.705 ;
        RECT 123.805 82.535 123.975 82.705 ;
        RECT 124.265 82.535 124.435 82.705 ;
        RECT 124.725 82.535 124.895 82.705 ;
        RECT 125.185 82.535 125.355 82.705 ;
        RECT 125.645 82.535 125.815 82.705 ;
        RECT 126.105 82.535 126.275 82.705 ;
        RECT 126.565 82.535 126.735 82.705 ;
        RECT 127.025 82.535 127.195 82.705 ;
        RECT 127.485 82.535 127.655 82.705 ;
        RECT 127.945 82.535 128.115 82.705 ;
        RECT 128.405 82.535 128.575 82.705 ;
        RECT 128.865 82.535 129.035 82.705 ;
        RECT 129.325 82.535 129.495 82.705 ;
        RECT 129.785 82.535 129.955 82.705 ;
        RECT 130.245 82.535 130.415 82.705 ;
        RECT 130.705 82.535 130.875 82.705 ;
        RECT 131.165 82.535 131.335 82.705 ;
        RECT 131.625 82.535 131.795 82.705 ;
        RECT 132.085 82.535 132.255 82.705 ;
        RECT 132.545 82.535 132.715 82.705 ;
        RECT 133.005 82.535 133.175 82.705 ;
        RECT 133.465 82.535 133.635 82.705 ;
        RECT 133.925 82.535 134.095 82.705 ;
        RECT 134.385 82.535 134.555 82.705 ;
        RECT 134.845 82.535 135.015 82.705 ;
        RECT 135.305 82.535 135.475 82.705 ;
        RECT 135.765 82.535 135.935 82.705 ;
        RECT 136.225 82.535 136.395 82.705 ;
        RECT 136.685 82.535 136.855 82.705 ;
        RECT 137.145 82.535 137.315 82.705 ;
        RECT 137.605 82.535 137.775 82.705 ;
        RECT 138.065 82.535 138.235 82.705 ;
        RECT 138.525 82.535 138.695 82.705 ;
        RECT 138.985 82.535 139.155 82.705 ;
        RECT 50.665 79.815 50.835 79.985 ;
        RECT 51.125 79.815 51.295 79.985 ;
        RECT 51.585 79.815 51.755 79.985 ;
        RECT 52.045 79.815 52.215 79.985 ;
        RECT 52.505 79.815 52.675 79.985 ;
        RECT 52.965 79.815 53.135 79.985 ;
        RECT 53.425 79.815 53.595 79.985 ;
        RECT 53.885 79.815 54.055 79.985 ;
        RECT 54.345 79.815 54.515 79.985 ;
        RECT 54.805 79.815 54.975 79.985 ;
        RECT 55.265 79.815 55.435 79.985 ;
        RECT 55.725 79.815 55.895 79.985 ;
        RECT 56.185 79.815 56.355 79.985 ;
        RECT 56.645 79.815 56.815 79.985 ;
        RECT 57.105 79.815 57.275 79.985 ;
        RECT 57.565 79.815 57.735 79.985 ;
        RECT 58.025 79.815 58.195 79.985 ;
        RECT 58.485 79.815 58.655 79.985 ;
        RECT 58.945 79.815 59.115 79.985 ;
        RECT 59.405 79.815 59.575 79.985 ;
        RECT 59.865 79.815 60.035 79.985 ;
        RECT 60.325 79.815 60.495 79.985 ;
        RECT 60.785 79.815 60.955 79.985 ;
        RECT 61.245 79.815 61.415 79.985 ;
        RECT 61.705 79.815 61.875 79.985 ;
        RECT 62.165 79.815 62.335 79.985 ;
        RECT 62.625 79.815 62.795 79.985 ;
        RECT 63.085 79.815 63.255 79.985 ;
        RECT 63.545 79.815 63.715 79.985 ;
        RECT 64.005 79.815 64.175 79.985 ;
        RECT 64.465 79.815 64.635 79.985 ;
        RECT 64.925 79.815 65.095 79.985 ;
        RECT 65.385 79.815 65.555 79.985 ;
        RECT 65.845 79.815 66.015 79.985 ;
        RECT 66.305 79.815 66.475 79.985 ;
        RECT 66.765 79.815 66.935 79.985 ;
        RECT 67.225 79.815 67.395 79.985 ;
        RECT 67.685 79.815 67.855 79.985 ;
        RECT 68.145 79.815 68.315 79.985 ;
        RECT 68.605 79.815 68.775 79.985 ;
        RECT 69.065 79.815 69.235 79.985 ;
        RECT 69.525 79.815 69.695 79.985 ;
        RECT 69.985 79.815 70.155 79.985 ;
        RECT 70.445 79.815 70.615 79.985 ;
        RECT 70.905 79.815 71.075 79.985 ;
        RECT 71.365 79.815 71.535 79.985 ;
        RECT 71.825 79.815 71.995 79.985 ;
        RECT 72.285 79.815 72.455 79.985 ;
        RECT 72.745 79.815 72.915 79.985 ;
        RECT 73.205 79.815 73.375 79.985 ;
        RECT 73.665 79.815 73.835 79.985 ;
        RECT 74.125 79.815 74.295 79.985 ;
        RECT 74.585 79.815 74.755 79.985 ;
        RECT 75.045 79.815 75.215 79.985 ;
        RECT 75.505 79.815 75.675 79.985 ;
        RECT 75.965 79.815 76.135 79.985 ;
        RECT 76.425 79.815 76.595 79.985 ;
        RECT 76.885 79.815 77.055 79.985 ;
        RECT 77.345 79.815 77.515 79.985 ;
        RECT 77.805 79.815 77.975 79.985 ;
        RECT 78.265 79.815 78.435 79.985 ;
        RECT 78.725 79.815 78.895 79.985 ;
        RECT 79.185 79.815 79.355 79.985 ;
        RECT 79.645 79.815 79.815 79.985 ;
        RECT 80.105 79.815 80.275 79.985 ;
        RECT 80.565 79.815 80.735 79.985 ;
        RECT 81.025 79.815 81.195 79.985 ;
        RECT 81.485 79.815 81.655 79.985 ;
        RECT 81.945 79.815 82.115 79.985 ;
        RECT 82.405 79.815 82.575 79.985 ;
        RECT 82.865 79.815 83.035 79.985 ;
        RECT 83.325 79.815 83.495 79.985 ;
        RECT 83.785 79.815 83.955 79.985 ;
        RECT 84.245 79.815 84.415 79.985 ;
        RECT 84.705 79.815 84.875 79.985 ;
        RECT 85.165 79.815 85.335 79.985 ;
        RECT 85.625 79.815 85.795 79.985 ;
        RECT 86.085 79.815 86.255 79.985 ;
        RECT 86.545 79.815 86.715 79.985 ;
        RECT 87.005 79.815 87.175 79.985 ;
        RECT 87.465 79.815 87.635 79.985 ;
        RECT 87.925 79.815 88.095 79.985 ;
        RECT 88.385 79.815 88.555 79.985 ;
        RECT 88.845 79.815 89.015 79.985 ;
        RECT 89.305 79.815 89.475 79.985 ;
        RECT 89.765 79.815 89.935 79.985 ;
        RECT 90.225 79.815 90.395 79.985 ;
        RECT 90.685 79.815 90.855 79.985 ;
        RECT 91.145 79.815 91.315 79.985 ;
        RECT 91.605 79.815 91.775 79.985 ;
        RECT 92.065 79.815 92.235 79.985 ;
        RECT 92.525 79.815 92.695 79.985 ;
        RECT 92.985 79.815 93.155 79.985 ;
        RECT 93.445 79.815 93.615 79.985 ;
        RECT 93.905 79.815 94.075 79.985 ;
        RECT 94.365 79.815 94.535 79.985 ;
        RECT 94.825 79.815 94.995 79.985 ;
        RECT 95.285 79.815 95.455 79.985 ;
        RECT 95.745 79.815 95.915 79.985 ;
        RECT 96.205 79.815 96.375 79.985 ;
        RECT 96.665 79.815 96.835 79.985 ;
        RECT 97.125 79.815 97.295 79.985 ;
        RECT 97.585 79.815 97.755 79.985 ;
        RECT 98.045 79.815 98.215 79.985 ;
        RECT 98.505 79.815 98.675 79.985 ;
        RECT 98.965 79.815 99.135 79.985 ;
        RECT 99.425 79.815 99.595 79.985 ;
        RECT 99.885 79.815 100.055 79.985 ;
        RECT 100.345 79.815 100.515 79.985 ;
        RECT 100.805 79.815 100.975 79.985 ;
        RECT 101.265 79.815 101.435 79.985 ;
        RECT 101.725 79.815 101.895 79.985 ;
        RECT 102.185 79.815 102.355 79.985 ;
        RECT 102.645 79.815 102.815 79.985 ;
        RECT 103.105 79.815 103.275 79.985 ;
        RECT 103.565 79.815 103.735 79.985 ;
        RECT 104.025 79.815 104.195 79.985 ;
        RECT 104.485 79.815 104.655 79.985 ;
        RECT 104.945 79.815 105.115 79.985 ;
        RECT 105.405 79.815 105.575 79.985 ;
        RECT 105.865 79.815 106.035 79.985 ;
        RECT 106.325 79.815 106.495 79.985 ;
        RECT 106.785 79.815 106.955 79.985 ;
        RECT 107.245 79.815 107.415 79.985 ;
        RECT 107.705 79.815 107.875 79.985 ;
        RECT 108.165 79.815 108.335 79.985 ;
        RECT 108.625 79.815 108.795 79.985 ;
        RECT 109.085 79.815 109.255 79.985 ;
        RECT 109.545 79.815 109.715 79.985 ;
        RECT 110.005 79.815 110.175 79.985 ;
        RECT 110.465 79.815 110.635 79.985 ;
        RECT 110.925 79.815 111.095 79.985 ;
        RECT 111.385 79.815 111.555 79.985 ;
        RECT 111.845 79.815 112.015 79.985 ;
        RECT 112.305 79.815 112.475 79.985 ;
        RECT 112.765 79.815 112.935 79.985 ;
        RECT 113.225 79.815 113.395 79.985 ;
        RECT 113.685 79.815 113.855 79.985 ;
        RECT 114.145 79.815 114.315 79.985 ;
        RECT 114.605 79.815 114.775 79.985 ;
        RECT 115.065 79.815 115.235 79.985 ;
        RECT 115.525 79.815 115.695 79.985 ;
        RECT 115.985 79.815 116.155 79.985 ;
        RECT 116.445 79.815 116.615 79.985 ;
        RECT 116.905 79.815 117.075 79.985 ;
        RECT 117.365 79.815 117.535 79.985 ;
        RECT 117.825 79.815 117.995 79.985 ;
        RECT 118.285 79.815 118.455 79.985 ;
        RECT 118.745 79.815 118.915 79.985 ;
        RECT 119.205 79.815 119.375 79.985 ;
        RECT 119.665 79.815 119.835 79.985 ;
        RECT 120.125 79.815 120.295 79.985 ;
        RECT 120.585 79.815 120.755 79.985 ;
        RECT 121.045 79.815 121.215 79.985 ;
        RECT 121.505 79.815 121.675 79.985 ;
        RECT 121.965 79.815 122.135 79.985 ;
        RECT 122.425 79.815 122.595 79.985 ;
        RECT 122.885 79.815 123.055 79.985 ;
        RECT 123.345 79.815 123.515 79.985 ;
        RECT 123.805 79.815 123.975 79.985 ;
        RECT 124.265 79.815 124.435 79.985 ;
        RECT 124.725 79.815 124.895 79.985 ;
        RECT 125.185 79.815 125.355 79.985 ;
        RECT 125.645 79.815 125.815 79.985 ;
        RECT 126.105 79.815 126.275 79.985 ;
        RECT 126.565 79.815 126.735 79.985 ;
        RECT 127.025 79.815 127.195 79.985 ;
        RECT 127.485 79.815 127.655 79.985 ;
        RECT 127.945 79.815 128.115 79.985 ;
        RECT 128.405 79.815 128.575 79.985 ;
        RECT 128.865 79.815 129.035 79.985 ;
        RECT 129.325 79.815 129.495 79.985 ;
        RECT 129.785 79.815 129.955 79.985 ;
        RECT 130.245 79.815 130.415 79.985 ;
        RECT 130.705 79.815 130.875 79.985 ;
        RECT 131.165 79.815 131.335 79.985 ;
        RECT 131.625 79.815 131.795 79.985 ;
        RECT 132.085 79.815 132.255 79.985 ;
        RECT 132.545 79.815 132.715 79.985 ;
        RECT 133.005 79.815 133.175 79.985 ;
        RECT 133.465 79.815 133.635 79.985 ;
        RECT 133.925 79.815 134.095 79.985 ;
        RECT 134.385 79.815 134.555 79.985 ;
        RECT 134.845 79.815 135.015 79.985 ;
        RECT 135.305 79.815 135.475 79.985 ;
        RECT 135.765 79.815 135.935 79.985 ;
        RECT 136.225 79.815 136.395 79.985 ;
        RECT 136.685 79.815 136.855 79.985 ;
        RECT 137.145 79.815 137.315 79.985 ;
        RECT 137.605 79.815 137.775 79.985 ;
        RECT 138.065 79.815 138.235 79.985 ;
        RECT 138.525 79.815 138.695 79.985 ;
        RECT 138.985 79.815 139.155 79.985 ;
        RECT 50.665 77.095 50.835 77.265 ;
        RECT 51.125 77.095 51.295 77.265 ;
        RECT 51.585 77.095 51.755 77.265 ;
        RECT 52.045 77.095 52.215 77.265 ;
        RECT 52.505 77.095 52.675 77.265 ;
        RECT 52.965 77.095 53.135 77.265 ;
        RECT 53.425 77.095 53.595 77.265 ;
        RECT 53.885 77.095 54.055 77.265 ;
        RECT 54.345 77.095 54.515 77.265 ;
        RECT 54.805 77.095 54.975 77.265 ;
        RECT 55.265 77.095 55.435 77.265 ;
        RECT 55.725 77.095 55.895 77.265 ;
        RECT 56.185 77.095 56.355 77.265 ;
        RECT 56.645 77.095 56.815 77.265 ;
        RECT 57.105 77.095 57.275 77.265 ;
        RECT 57.565 77.095 57.735 77.265 ;
        RECT 58.025 77.095 58.195 77.265 ;
        RECT 58.485 77.095 58.655 77.265 ;
        RECT 58.945 77.095 59.115 77.265 ;
        RECT 59.405 77.095 59.575 77.265 ;
        RECT 59.865 77.095 60.035 77.265 ;
        RECT 60.325 77.095 60.495 77.265 ;
        RECT 60.785 77.095 60.955 77.265 ;
        RECT 61.245 77.095 61.415 77.265 ;
        RECT 61.705 77.095 61.875 77.265 ;
        RECT 62.165 77.095 62.335 77.265 ;
        RECT 62.625 77.095 62.795 77.265 ;
        RECT 63.085 77.095 63.255 77.265 ;
        RECT 63.545 77.095 63.715 77.265 ;
        RECT 64.005 77.095 64.175 77.265 ;
        RECT 64.465 77.095 64.635 77.265 ;
        RECT 64.925 77.095 65.095 77.265 ;
        RECT 65.385 77.095 65.555 77.265 ;
        RECT 65.845 77.095 66.015 77.265 ;
        RECT 66.305 77.095 66.475 77.265 ;
        RECT 66.765 77.095 66.935 77.265 ;
        RECT 67.225 77.095 67.395 77.265 ;
        RECT 67.685 77.095 67.855 77.265 ;
        RECT 68.145 77.095 68.315 77.265 ;
        RECT 68.605 77.095 68.775 77.265 ;
        RECT 69.065 77.095 69.235 77.265 ;
        RECT 69.525 77.095 69.695 77.265 ;
        RECT 69.985 77.095 70.155 77.265 ;
        RECT 70.445 77.095 70.615 77.265 ;
        RECT 70.905 77.095 71.075 77.265 ;
        RECT 71.365 77.095 71.535 77.265 ;
        RECT 71.825 77.095 71.995 77.265 ;
        RECT 72.285 77.095 72.455 77.265 ;
        RECT 72.745 77.095 72.915 77.265 ;
        RECT 73.205 77.095 73.375 77.265 ;
        RECT 73.665 77.095 73.835 77.265 ;
        RECT 74.125 77.095 74.295 77.265 ;
        RECT 74.585 77.095 74.755 77.265 ;
        RECT 75.045 77.095 75.215 77.265 ;
        RECT 75.505 77.095 75.675 77.265 ;
        RECT 75.965 77.095 76.135 77.265 ;
        RECT 76.425 77.095 76.595 77.265 ;
        RECT 76.885 77.095 77.055 77.265 ;
        RECT 77.345 77.095 77.515 77.265 ;
        RECT 77.805 77.095 77.975 77.265 ;
        RECT 78.265 77.095 78.435 77.265 ;
        RECT 78.725 77.095 78.895 77.265 ;
        RECT 79.185 77.095 79.355 77.265 ;
        RECT 79.645 77.095 79.815 77.265 ;
        RECT 80.105 77.095 80.275 77.265 ;
        RECT 80.565 77.095 80.735 77.265 ;
        RECT 81.025 77.095 81.195 77.265 ;
        RECT 81.485 77.095 81.655 77.265 ;
        RECT 81.945 77.095 82.115 77.265 ;
        RECT 82.405 77.095 82.575 77.265 ;
        RECT 82.865 77.095 83.035 77.265 ;
        RECT 83.325 77.095 83.495 77.265 ;
        RECT 83.785 77.095 83.955 77.265 ;
        RECT 84.245 77.095 84.415 77.265 ;
        RECT 84.705 77.095 84.875 77.265 ;
        RECT 85.165 77.095 85.335 77.265 ;
        RECT 85.625 77.095 85.795 77.265 ;
        RECT 86.085 77.095 86.255 77.265 ;
        RECT 86.545 77.095 86.715 77.265 ;
        RECT 87.005 77.095 87.175 77.265 ;
        RECT 87.465 77.095 87.635 77.265 ;
        RECT 87.925 77.095 88.095 77.265 ;
        RECT 88.385 77.095 88.555 77.265 ;
        RECT 88.845 77.095 89.015 77.265 ;
        RECT 89.305 77.095 89.475 77.265 ;
        RECT 89.765 77.095 89.935 77.265 ;
        RECT 90.225 77.095 90.395 77.265 ;
        RECT 90.685 77.095 90.855 77.265 ;
        RECT 91.145 77.095 91.315 77.265 ;
        RECT 91.605 77.095 91.775 77.265 ;
        RECT 92.065 77.095 92.235 77.265 ;
        RECT 92.525 77.095 92.695 77.265 ;
        RECT 92.985 77.095 93.155 77.265 ;
        RECT 93.445 77.095 93.615 77.265 ;
        RECT 93.905 77.095 94.075 77.265 ;
        RECT 94.365 77.095 94.535 77.265 ;
        RECT 94.825 77.095 94.995 77.265 ;
        RECT 95.285 77.095 95.455 77.265 ;
        RECT 95.745 77.095 95.915 77.265 ;
        RECT 96.205 77.095 96.375 77.265 ;
        RECT 96.665 77.095 96.835 77.265 ;
        RECT 97.125 77.095 97.295 77.265 ;
        RECT 97.585 77.095 97.755 77.265 ;
        RECT 98.045 77.095 98.215 77.265 ;
        RECT 98.505 77.095 98.675 77.265 ;
        RECT 98.965 77.095 99.135 77.265 ;
        RECT 99.425 77.095 99.595 77.265 ;
        RECT 99.885 77.095 100.055 77.265 ;
        RECT 100.345 77.095 100.515 77.265 ;
        RECT 100.805 77.095 100.975 77.265 ;
        RECT 101.265 77.095 101.435 77.265 ;
        RECT 101.725 77.095 101.895 77.265 ;
        RECT 102.185 77.095 102.355 77.265 ;
        RECT 102.645 77.095 102.815 77.265 ;
        RECT 103.105 77.095 103.275 77.265 ;
        RECT 103.565 77.095 103.735 77.265 ;
        RECT 104.025 77.095 104.195 77.265 ;
        RECT 104.485 77.095 104.655 77.265 ;
        RECT 104.945 77.095 105.115 77.265 ;
        RECT 105.405 77.095 105.575 77.265 ;
        RECT 105.865 77.095 106.035 77.265 ;
        RECT 106.325 77.095 106.495 77.265 ;
        RECT 106.785 77.095 106.955 77.265 ;
        RECT 107.245 77.095 107.415 77.265 ;
        RECT 107.705 77.095 107.875 77.265 ;
        RECT 108.165 77.095 108.335 77.265 ;
        RECT 108.625 77.095 108.795 77.265 ;
        RECT 109.085 77.095 109.255 77.265 ;
        RECT 109.545 77.095 109.715 77.265 ;
        RECT 110.005 77.095 110.175 77.265 ;
        RECT 110.465 77.095 110.635 77.265 ;
        RECT 110.925 77.095 111.095 77.265 ;
        RECT 111.385 77.095 111.555 77.265 ;
        RECT 111.845 77.095 112.015 77.265 ;
        RECT 112.305 77.095 112.475 77.265 ;
        RECT 112.765 77.095 112.935 77.265 ;
        RECT 113.225 77.095 113.395 77.265 ;
        RECT 113.685 77.095 113.855 77.265 ;
        RECT 114.145 77.095 114.315 77.265 ;
        RECT 114.605 77.095 114.775 77.265 ;
        RECT 115.065 77.095 115.235 77.265 ;
        RECT 115.525 77.095 115.695 77.265 ;
        RECT 115.985 77.095 116.155 77.265 ;
        RECT 116.445 77.095 116.615 77.265 ;
        RECT 116.905 77.095 117.075 77.265 ;
        RECT 117.365 77.095 117.535 77.265 ;
        RECT 117.825 77.095 117.995 77.265 ;
        RECT 118.285 77.095 118.455 77.265 ;
        RECT 118.745 77.095 118.915 77.265 ;
        RECT 119.205 77.095 119.375 77.265 ;
        RECT 119.665 77.095 119.835 77.265 ;
        RECT 120.125 77.095 120.295 77.265 ;
        RECT 120.585 77.095 120.755 77.265 ;
        RECT 121.045 77.095 121.215 77.265 ;
        RECT 121.505 77.095 121.675 77.265 ;
        RECT 121.965 77.095 122.135 77.265 ;
        RECT 122.425 77.095 122.595 77.265 ;
        RECT 122.885 77.095 123.055 77.265 ;
        RECT 123.345 77.095 123.515 77.265 ;
        RECT 123.805 77.095 123.975 77.265 ;
        RECT 124.265 77.095 124.435 77.265 ;
        RECT 124.725 77.095 124.895 77.265 ;
        RECT 125.185 77.095 125.355 77.265 ;
        RECT 125.645 77.095 125.815 77.265 ;
        RECT 126.105 77.095 126.275 77.265 ;
        RECT 126.565 77.095 126.735 77.265 ;
        RECT 127.025 77.095 127.195 77.265 ;
        RECT 127.485 77.095 127.655 77.265 ;
        RECT 127.945 77.095 128.115 77.265 ;
        RECT 128.405 77.095 128.575 77.265 ;
        RECT 128.865 77.095 129.035 77.265 ;
        RECT 129.325 77.095 129.495 77.265 ;
        RECT 129.785 77.095 129.955 77.265 ;
        RECT 130.245 77.095 130.415 77.265 ;
        RECT 130.705 77.095 130.875 77.265 ;
        RECT 131.165 77.095 131.335 77.265 ;
        RECT 131.625 77.095 131.795 77.265 ;
        RECT 132.085 77.095 132.255 77.265 ;
        RECT 132.545 77.095 132.715 77.265 ;
        RECT 133.005 77.095 133.175 77.265 ;
        RECT 133.465 77.095 133.635 77.265 ;
        RECT 133.925 77.095 134.095 77.265 ;
        RECT 134.385 77.095 134.555 77.265 ;
        RECT 134.845 77.095 135.015 77.265 ;
        RECT 135.305 77.095 135.475 77.265 ;
        RECT 135.765 77.095 135.935 77.265 ;
        RECT 136.225 77.095 136.395 77.265 ;
        RECT 136.685 77.095 136.855 77.265 ;
        RECT 137.145 77.095 137.315 77.265 ;
        RECT 137.605 77.095 137.775 77.265 ;
        RECT 138.065 77.095 138.235 77.265 ;
        RECT 138.525 77.095 138.695 77.265 ;
        RECT 138.985 77.095 139.155 77.265 ;
        RECT 50.665 74.375 50.835 74.545 ;
        RECT 51.125 74.375 51.295 74.545 ;
        RECT 51.585 74.375 51.755 74.545 ;
        RECT 52.045 74.375 52.215 74.545 ;
        RECT 52.505 74.375 52.675 74.545 ;
        RECT 52.965 74.375 53.135 74.545 ;
        RECT 53.425 74.375 53.595 74.545 ;
        RECT 53.885 74.375 54.055 74.545 ;
        RECT 54.345 74.375 54.515 74.545 ;
        RECT 54.805 74.375 54.975 74.545 ;
        RECT 55.265 74.375 55.435 74.545 ;
        RECT 55.725 74.375 55.895 74.545 ;
        RECT 56.185 74.375 56.355 74.545 ;
        RECT 56.645 74.375 56.815 74.545 ;
        RECT 57.105 74.375 57.275 74.545 ;
        RECT 57.565 74.375 57.735 74.545 ;
        RECT 58.025 74.375 58.195 74.545 ;
        RECT 58.485 74.375 58.655 74.545 ;
        RECT 58.945 74.375 59.115 74.545 ;
        RECT 59.405 74.375 59.575 74.545 ;
        RECT 59.865 74.375 60.035 74.545 ;
        RECT 60.325 74.375 60.495 74.545 ;
        RECT 60.785 74.375 60.955 74.545 ;
        RECT 61.245 74.375 61.415 74.545 ;
        RECT 61.705 74.375 61.875 74.545 ;
        RECT 62.165 74.375 62.335 74.545 ;
        RECT 62.625 74.375 62.795 74.545 ;
        RECT 63.085 74.375 63.255 74.545 ;
        RECT 63.545 74.375 63.715 74.545 ;
        RECT 64.005 74.375 64.175 74.545 ;
        RECT 64.465 74.375 64.635 74.545 ;
        RECT 64.925 74.375 65.095 74.545 ;
        RECT 65.385 74.375 65.555 74.545 ;
        RECT 65.845 74.375 66.015 74.545 ;
        RECT 66.305 74.375 66.475 74.545 ;
        RECT 66.765 74.375 66.935 74.545 ;
        RECT 67.225 74.375 67.395 74.545 ;
        RECT 67.685 74.375 67.855 74.545 ;
        RECT 68.145 74.375 68.315 74.545 ;
        RECT 68.605 74.375 68.775 74.545 ;
        RECT 69.065 74.375 69.235 74.545 ;
        RECT 69.525 74.375 69.695 74.545 ;
        RECT 69.985 74.375 70.155 74.545 ;
        RECT 70.445 74.375 70.615 74.545 ;
        RECT 70.905 74.375 71.075 74.545 ;
        RECT 71.365 74.375 71.535 74.545 ;
        RECT 71.825 74.375 71.995 74.545 ;
        RECT 72.285 74.375 72.455 74.545 ;
        RECT 72.745 74.375 72.915 74.545 ;
        RECT 73.205 74.375 73.375 74.545 ;
        RECT 73.665 74.375 73.835 74.545 ;
        RECT 74.125 74.375 74.295 74.545 ;
        RECT 74.585 74.375 74.755 74.545 ;
        RECT 75.045 74.375 75.215 74.545 ;
        RECT 75.505 74.375 75.675 74.545 ;
        RECT 75.965 74.375 76.135 74.545 ;
        RECT 76.425 74.375 76.595 74.545 ;
        RECT 76.885 74.375 77.055 74.545 ;
        RECT 77.345 74.375 77.515 74.545 ;
        RECT 77.805 74.375 77.975 74.545 ;
        RECT 78.265 74.375 78.435 74.545 ;
        RECT 78.725 74.375 78.895 74.545 ;
        RECT 79.185 74.375 79.355 74.545 ;
        RECT 79.645 74.375 79.815 74.545 ;
        RECT 80.105 74.375 80.275 74.545 ;
        RECT 80.565 74.375 80.735 74.545 ;
        RECT 81.025 74.375 81.195 74.545 ;
        RECT 81.485 74.375 81.655 74.545 ;
        RECT 81.945 74.375 82.115 74.545 ;
        RECT 82.405 74.375 82.575 74.545 ;
        RECT 82.865 74.375 83.035 74.545 ;
        RECT 83.325 74.375 83.495 74.545 ;
        RECT 83.785 74.375 83.955 74.545 ;
        RECT 84.245 74.375 84.415 74.545 ;
        RECT 84.705 74.375 84.875 74.545 ;
        RECT 85.165 74.375 85.335 74.545 ;
        RECT 85.625 74.375 85.795 74.545 ;
        RECT 86.085 74.375 86.255 74.545 ;
        RECT 86.545 74.375 86.715 74.545 ;
        RECT 87.005 74.375 87.175 74.545 ;
        RECT 87.465 74.375 87.635 74.545 ;
        RECT 87.925 74.375 88.095 74.545 ;
        RECT 88.385 74.375 88.555 74.545 ;
        RECT 88.845 74.375 89.015 74.545 ;
        RECT 89.305 74.375 89.475 74.545 ;
        RECT 89.765 74.375 89.935 74.545 ;
        RECT 90.225 74.375 90.395 74.545 ;
        RECT 90.685 74.375 90.855 74.545 ;
        RECT 91.145 74.375 91.315 74.545 ;
        RECT 91.605 74.375 91.775 74.545 ;
        RECT 92.065 74.375 92.235 74.545 ;
        RECT 92.525 74.375 92.695 74.545 ;
        RECT 92.985 74.375 93.155 74.545 ;
        RECT 93.445 74.375 93.615 74.545 ;
        RECT 93.905 74.375 94.075 74.545 ;
        RECT 94.365 74.375 94.535 74.545 ;
        RECT 94.825 74.375 94.995 74.545 ;
        RECT 95.285 74.375 95.455 74.545 ;
        RECT 95.745 74.375 95.915 74.545 ;
        RECT 96.205 74.375 96.375 74.545 ;
        RECT 96.665 74.375 96.835 74.545 ;
        RECT 97.125 74.375 97.295 74.545 ;
        RECT 97.585 74.375 97.755 74.545 ;
        RECT 98.045 74.375 98.215 74.545 ;
        RECT 98.505 74.375 98.675 74.545 ;
        RECT 98.965 74.375 99.135 74.545 ;
        RECT 99.425 74.375 99.595 74.545 ;
        RECT 99.885 74.375 100.055 74.545 ;
        RECT 100.345 74.375 100.515 74.545 ;
        RECT 100.805 74.375 100.975 74.545 ;
        RECT 101.265 74.375 101.435 74.545 ;
        RECT 101.725 74.375 101.895 74.545 ;
        RECT 102.185 74.375 102.355 74.545 ;
        RECT 102.645 74.375 102.815 74.545 ;
        RECT 103.105 74.375 103.275 74.545 ;
        RECT 103.565 74.375 103.735 74.545 ;
        RECT 104.025 74.375 104.195 74.545 ;
        RECT 104.485 74.375 104.655 74.545 ;
        RECT 104.945 74.375 105.115 74.545 ;
        RECT 105.405 74.375 105.575 74.545 ;
        RECT 105.865 74.375 106.035 74.545 ;
        RECT 106.325 74.375 106.495 74.545 ;
        RECT 106.785 74.375 106.955 74.545 ;
        RECT 107.245 74.375 107.415 74.545 ;
        RECT 107.705 74.375 107.875 74.545 ;
        RECT 108.165 74.375 108.335 74.545 ;
        RECT 108.625 74.375 108.795 74.545 ;
        RECT 109.085 74.375 109.255 74.545 ;
        RECT 109.545 74.375 109.715 74.545 ;
        RECT 110.005 74.375 110.175 74.545 ;
        RECT 110.465 74.375 110.635 74.545 ;
        RECT 110.925 74.375 111.095 74.545 ;
        RECT 111.385 74.375 111.555 74.545 ;
        RECT 111.845 74.375 112.015 74.545 ;
        RECT 112.305 74.375 112.475 74.545 ;
        RECT 112.765 74.375 112.935 74.545 ;
        RECT 113.225 74.375 113.395 74.545 ;
        RECT 113.685 74.375 113.855 74.545 ;
        RECT 114.145 74.375 114.315 74.545 ;
        RECT 114.605 74.375 114.775 74.545 ;
        RECT 115.065 74.375 115.235 74.545 ;
        RECT 115.525 74.375 115.695 74.545 ;
        RECT 115.985 74.375 116.155 74.545 ;
        RECT 116.445 74.375 116.615 74.545 ;
        RECT 116.905 74.375 117.075 74.545 ;
        RECT 117.365 74.375 117.535 74.545 ;
        RECT 117.825 74.375 117.995 74.545 ;
        RECT 118.285 74.375 118.455 74.545 ;
        RECT 118.745 74.375 118.915 74.545 ;
        RECT 119.205 74.375 119.375 74.545 ;
        RECT 119.665 74.375 119.835 74.545 ;
        RECT 120.125 74.375 120.295 74.545 ;
        RECT 120.585 74.375 120.755 74.545 ;
        RECT 121.045 74.375 121.215 74.545 ;
        RECT 121.505 74.375 121.675 74.545 ;
        RECT 121.965 74.375 122.135 74.545 ;
        RECT 122.425 74.375 122.595 74.545 ;
        RECT 122.885 74.375 123.055 74.545 ;
        RECT 123.345 74.375 123.515 74.545 ;
        RECT 123.805 74.375 123.975 74.545 ;
        RECT 124.265 74.375 124.435 74.545 ;
        RECT 124.725 74.375 124.895 74.545 ;
        RECT 125.185 74.375 125.355 74.545 ;
        RECT 125.645 74.375 125.815 74.545 ;
        RECT 126.105 74.375 126.275 74.545 ;
        RECT 126.565 74.375 126.735 74.545 ;
        RECT 127.025 74.375 127.195 74.545 ;
        RECT 127.485 74.375 127.655 74.545 ;
        RECT 127.945 74.375 128.115 74.545 ;
        RECT 128.405 74.375 128.575 74.545 ;
        RECT 128.865 74.375 129.035 74.545 ;
        RECT 129.325 74.375 129.495 74.545 ;
        RECT 129.785 74.375 129.955 74.545 ;
        RECT 130.245 74.375 130.415 74.545 ;
        RECT 130.705 74.375 130.875 74.545 ;
        RECT 131.165 74.375 131.335 74.545 ;
        RECT 131.625 74.375 131.795 74.545 ;
        RECT 132.085 74.375 132.255 74.545 ;
        RECT 132.545 74.375 132.715 74.545 ;
        RECT 133.005 74.375 133.175 74.545 ;
        RECT 133.465 74.375 133.635 74.545 ;
        RECT 133.925 74.375 134.095 74.545 ;
        RECT 134.385 74.375 134.555 74.545 ;
        RECT 134.845 74.375 135.015 74.545 ;
        RECT 135.305 74.375 135.475 74.545 ;
        RECT 135.765 74.375 135.935 74.545 ;
        RECT 136.225 74.375 136.395 74.545 ;
        RECT 136.685 74.375 136.855 74.545 ;
        RECT 137.145 74.375 137.315 74.545 ;
        RECT 137.605 74.375 137.775 74.545 ;
        RECT 138.065 74.375 138.235 74.545 ;
        RECT 138.525 74.375 138.695 74.545 ;
        RECT 138.985 74.375 139.155 74.545 ;
        RECT 50.665 71.655 50.835 71.825 ;
        RECT 51.125 71.655 51.295 71.825 ;
        RECT 51.585 71.655 51.755 71.825 ;
        RECT 52.045 71.655 52.215 71.825 ;
        RECT 52.505 71.655 52.675 71.825 ;
        RECT 52.965 71.655 53.135 71.825 ;
        RECT 53.425 71.655 53.595 71.825 ;
        RECT 53.885 71.655 54.055 71.825 ;
        RECT 54.345 71.655 54.515 71.825 ;
        RECT 54.805 71.655 54.975 71.825 ;
        RECT 55.265 71.655 55.435 71.825 ;
        RECT 55.725 71.655 55.895 71.825 ;
        RECT 56.185 71.655 56.355 71.825 ;
        RECT 56.645 71.655 56.815 71.825 ;
        RECT 57.105 71.655 57.275 71.825 ;
        RECT 57.565 71.655 57.735 71.825 ;
        RECT 58.025 71.655 58.195 71.825 ;
        RECT 58.485 71.655 58.655 71.825 ;
        RECT 58.945 71.655 59.115 71.825 ;
        RECT 59.405 71.655 59.575 71.825 ;
        RECT 59.865 71.655 60.035 71.825 ;
        RECT 60.325 71.655 60.495 71.825 ;
        RECT 60.785 71.655 60.955 71.825 ;
        RECT 61.245 71.655 61.415 71.825 ;
        RECT 61.705 71.655 61.875 71.825 ;
        RECT 62.165 71.655 62.335 71.825 ;
        RECT 62.625 71.655 62.795 71.825 ;
        RECT 63.085 71.655 63.255 71.825 ;
        RECT 63.545 71.655 63.715 71.825 ;
        RECT 64.005 71.655 64.175 71.825 ;
        RECT 64.465 71.655 64.635 71.825 ;
        RECT 64.925 71.655 65.095 71.825 ;
        RECT 65.385 71.655 65.555 71.825 ;
        RECT 65.845 71.655 66.015 71.825 ;
        RECT 66.305 71.655 66.475 71.825 ;
        RECT 66.765 71.655 66.935 71.825 ;
        RECT 67.225 71.655 67.395 71.825 ;
        RECT 67.685 71.655 67.855 71.825 ;
        RECT 68.145 71.655 68.315 71.825 ;
        RECT 68.605 71.655 68.775 71.825 ;
        RECT 69.065 71.655 69.235 71.825 ;
        RECT 69.525 71.655 69.695 71.825 ;
        RECT 69.985 71.655 70.155 71.825 ;
        RECT 70.445 71.655 70.615 71.825 ;
        RECT 70.905 71.655 71.075 71.825 ;
        RECT 71.365 71.655 71.535 71.825 ;
        RECT 71.825 71.655 71.995 71.825 ;
        RECT 72.285 71.655 72.455 71.825 ;
        RECT 72.745 71.655 72.915 71.825 ;
        RECT 73.205 71.655 73.375 71.825 ;
        RECT 73.665 71.655 73.835 71.825 ;
        RECT 74.125 71.655 74.295 71.825 ;
        RECT 74.585 71.655 74.755 71.825 ;
        RECT 75.045 71.655 75.215 71.825 ;
        RECT 75.505 71.655 75.675 71.825 ;
        RECT 75.965 71.655 76.135 71.825 ;
        RECT 76.425 71.655 76.595 71.825 ;
        RECT 76.885 71.655 77.055 71.825 ;
        RECT 77.345 71.655 77.515 71.825 ;
        RECT 77.805 71.655 77.975 71.825 ;
        RECT 78.265 71.655 78.435 71.825 ;
        RECT 78.725 71.655 78.895 71.825 ;
        RECT 79.185 71.655 79.355 71.825 ;
        RECT 79.645 71.655 79.815 71.825 ;
        RECT 80.105 71.655 80.275 71.825 ;
        RECT 80.565 71.655 80.735 71.825 ;
        RECT 81.025 71.655 81.195 71.825 ;
        RECT 81.485 71.655 81.655 71.825 ;
        RECT 81.945 71.655 82.115 71.825 ;
        RECT 82.405 71.655 82.575 71.825 ;
        RECT 82.865 71.655 83.035 71.825 ;
        RECT 83.325 71.655 83.495 71.825 ;
        RECT 83.785 71.655 83.955 71.825 ;
        RECT 84.245 71.655 84.415 71.825 ;
        RECT 84.705 71.655 84.875 71.825 ;
        RECT 85.165 71.655 85.335 71.825 ;
        RECT 85.625 71.655 85.795 71.825 ;
        RECT 86.085 71.655 86.255 71.825 ;
        RECT 86.545 71.655 86.715 71.825 ;
        RECT 87.005 71.655 87.175 71.825 ;
        RECT 87.465 71.655 87.635 71.825 ;
        RECT 87.925 71.655 88.095 71.825 ;
        RECT 88.385 71.655 88.555 71.825 ;
        RECT 88.845 71.655 89.015 71.825 ;
        RECT 89.305 71.655 89.475 71.825 ;
        RECT 89.765 71.655 89.935 71.825 ;
        RECT 90.225 71.655 90.395 71.825 ;
        RECT 90.685 71.655 90.855 71.825 ;
        RECT 91.145 71.655 91.315 71.825 ;
        RECT 91.605 71.655 91.775 71.825 ;
        RECT 92.065 71.655 92.235 71.825 ;
        RECT 92.525 71.655 92.695 71.825 ;
        RECT 92.985 71.655 93.155 71.825 ;
        RECT 93.445 71.655 93.615 71.825 ;
        RECT 93.905 71.655 94.075 71.825 ;
        RECT 94.365 71.655 94.535 71.825 ;
        RECT 94.825 71.655 94.995 71.825 ;
        RECT 95.285 71.655 95.455 71.825 ;
        RECT 95.745 71.655 95.915 71.825 ;
        RECT 96.205 71.655 96.375 71.825 ;
        RECT 96.665 71.655 96.835 71.825 ;
        RECT 97.125 71.655 97.295 71.825 ;
        RECT 97.585 71.655 97.755 71.825 ;
        RECT 98.045 71.655 98.215 71.825 ;
        RECT 98.505 71.655 98.675 71.825 ;
        RECT 98.965 71.655 99.135 71.825 ;
        RECT 99.425 71.655 99.595 71.825 ;
        RECT 99.885 71.655 100.055 71.825 ;
        RECT 100.345 71.655 100.515 71.825 ;
        RECT 100.805 71.655 100.975 71.825 ;
        RECT 101.265 71.655 101.435 71.825 ;
        RECT 101.725 71.655 101.895 71.825 ;
        RECT 102.185 71.655 102.355 71.825 ;
        RECT 102.645 71.655 102.815 71.825 ;
        RECT 103.105 71.655 103.275 71.825 ;
        RECT 103.565 71.655 103.735 71.825 ;
        RECT 104.025 71.655 104.195 71.825 ;
        RECT 104.485 71.655 104.655 71.825 ;
        RECT 104.945 71.655 105.115 71.825 ;
        RECT 105.405 71.655 105.575 71.825 ;
        RECT 105.865 71.655 106.035 71.825 ;
        RECT 106.325 71.655 106.495 71.825 ;
        RECT 106.785 71.655 106.955 71.825 ;
        RECT 107.245 71.655 107.415 71.825 ;
        RECT 107.705 71.655 107.875 71.825 ;
        RECT 108.165 71.655 108.335 71.825 ;
        RECT 108.625 71.655 108.795 71.825 ;
        RECT 109.085 71.655 109.255 71.825 ;
        RECT 109.545 71.655 109.715 71.825 ;
        RECT 110.005 71.655 110.175 71.825 ;
        RECT 110.465 71.655 110.635 71.825 ;
        RECT 110.925 71.655 111.095 71.825 ;
        RECT 111.385 71.655 111.555 71.825 ;
        RECT 111.845 71.655 112.015 71.825 ;
        RECT 112.305 71.655 112.475 71.825 ;
        RECT 112.765 71.655 112.935 71.825 ;
        RECT 113.225 71.655 113.395 71.825 ;
        RECT 113.685 71.655 113.855 71.825 ;
        RECT 114.145 71.655 114.315 71.825 ;
        RECT 114.605 71.655 114.775 71.825 ;
        RECT 115.065 71.655 115.235 71.825 ;
        RECT 115.525 71.655 115.695 71.825 ;
        RECT 115.985 71.655 116.155 71.825 ;
        RECT 116.445 71.655 116.615 71.825 ;
        RECT 116.905 71.655 117.075 71.825 ;
        RECT 117.365 71.655 117.535 71.825 ;
        RECT 117.825 71.655 117.995 71.825 ;
        RECT 118.285 71.655 118.455 71.825 ;
        RECT 118.745 71.655 118.915 71.825 ;
        RECT 119.205 71.655 119.375 71.825 ;
        RECT 119.665 71.655 119.835 71.825 ;
        RECT 120.125 71.655 120.295 71.825 ;
        RECT 120.585 71.655 120.755 71.825 ;
        RECT 121.045 71.655 121.215 71.825 ;
        RECT 121.505 71.655 121.675 71.825 ;
        RECT 121.965 71.655 122.135 71.825 ;
        RECT 122.425 71.655 122.595 71.825 ;
        RECT 122.885 71.655 123.055 71.825 ;
        RECT 123.345 71.655 123.515 71.825 ;
        RECT 123.805 71.655 123.975 71.825 ;
        RECT 124.265 71.655 124.435 71.825 ;
        RECT 124.725 71.655 124.895 71.825 ;
        RECT 125.185 71.655 125.355 71.825 ;
        RECT 125.645 71.655 125.815 71.825 ;
        RECT 126.105 71.655 126.275 71.825 ;
        RECT 126.565 71.655 126.735 71.825 ;
        RECT 127.025 71.655 127.195 71.825 ;
        RECT 127.485 71.655 127.655 71.825 ;
        RECT 127.945 71.655 128.115 71.825 ;
        RECT 128.405 71.655 128.575 71.825 ;
        RECT 128.865 71.655 129.035 71.825 ;
        RECT 129.325 71.655 129.495 71.825 ;
        RECT 129.785 71.655 129.955 71.825 ;
        RECT 130.245 71.655 130.415 71.825 ;
        RECT 130.705 71.655 130.875 71.825 ;
        RECT 131.165 71.655 131.335 71.825 ;
        RECT 131.625 71.655 131.795 71.825 ;
        RECT 132.085 71.655 132.255 71.825 ;
        RECT 132.545 71.655 132.715 71.825 ;
        RECT 133.005 71.655 133.175 71.825 ;
        RECT 133.465 71.655 133.635 71.825 ;
        RECT 133.925 71.655 134.095 71.825 ;
        RECT 134.385 71.655 134.555 71.825 ;
        RECT 134.845 71.655 135.015 71.825 ;
        RECT 135.305 71.655 135.475 71.825 ;
        RECT 135.765 71.655 135.935 71.825 ;
        RECT 136.225 71.655 136.395 71.825 ;
        RECT 136.685 71.655 136.855 71.825 ;
        RECT 137.145 71.655 137.315 71.825 ;
        RECT 137.605 71.655 137.775 71.825 ;
        RECT 138.065 71.655 138.235 71.825 ;
        RECT 138.525 71.655 138.695 71.825 ;
        RECT 138.985 71.655 139.155 71.825 ;
        RECT 50.665 68.935 50.835 69.105 ;
        RECT 51.125 68.935 51.295 69.105 ;
        RECT 51.585 68.935 51.755 69.105 ;
        RECT 52.045 68.935 52.215 69.105 ;
        RECT 52.505 68.935 52.675 69.105 ;
        RECT 52.965 68.935 53.135 69.105 ;
        RECT 53.425 68.935 53.595 69.105 ;
        RECT 53.885 68.935 54.055 69.105 ;
        RECT 54.345 68.935 54.515 69.105 ;
        RECT 54.805 68.935 54.975 69.105 ;
        RECT 55.265 68.935 55.435 69.105 ;
        RECT 55.725 68.935 55.895 69.105 ;
        RECT 56.185 68.935 56.355 69.105 ;
        RECT 56.645 68.935 56.815 69.105 ;
        RECT 57.105 68.935 57.275 69.105 ;
        RECT 57.565 68.935 57.735 69.105 ;
        RECT 58.025 68.935 58.195 69.105 ;
        RECT 58.485 68.935 58.655 69.105 ;
        RECT 58.945 68.935 59.115 69.105 ;
        RECT 59.405 68.935 59.575 69.105 ;
        RECT 59.865 68.935 60.035 69.105 ;
        RECT 60.325 68.935 60.495 69.105 ;
        RECT 60.785 68.935 60.955 69.105 ;
        RECT 61.245 68.935 61.415 69.105 ;
        RECT 61.705 68.935 61.875 69.105 ;
        RECT 62.165 68.935 62.335 69.105 ;
        RECT 62.625 68.935 62.795 69.105 ;
        RECT 63.085 68.935 63.255 69.105 ;
        RECT 63.545 68.935 63.715 69.105 ;
        RECT 64.005 68.935 64.175 69.105 ;
        RECT 64.465 68.935 64.635 69.105 ;
        RECT 64.925 68.935 65.095 69.105 ;
        RECT 65.385 68.935 65.555 69.105 ;
        RECT 65.845 68.935 66.015 69.105 ;
        RECT 66.305 68.935 66.475 69.105 ;
        RECT 66.765 68.935 66.935 69.105 ;
        RECT 67.225 68.935 67.395 69.105 ;
        RECT 67.685 68.935 67.855 69.105 ;
        RECT 68.145 68.935 68.315 69.105 ;
        RECT 68.605 68.935 68.775 69.105 ;
        RECT 69.065 68.935 69.235 69.105 ;
        RECT 69.525 68.935 69.695 69.105 ;
        RECT 69.985 68.935 70.155 69.105 ;
        RECT 70.445 68.935 70.615 69.105 ;
        RECT 70.905 68.935 71.075 69.105 ;
        RECT 71.365 68.935 71.535 69.105 ;
        RECT 71.825 68.935 71.995 69.105 ;
        RECT 72.285 68.935 72.455 69.105 ;
        RECT 72.745 68.935 72.915 69.105 ;
        RECT 73.205 68.935 73.375 69.105 ;
        RECT 73.665 68.935 73.835 69.105 ;
        RECT 74.125 68.935 74.295 69.105 ;
        RECT 74.585 68.935 74.755 69.105 ;
        RECT 75.045 68.935 75.215 69.105 ;
        RECT 75.505 68.935 75.675 69.105 ;
        RECT 75.965 68.935 76.135 69.105 ;
        RECT 76.425 68.935 76.595 69.105 ;
        RECT 76.885 68.935 77.055 69.105 ;
        RECT 77.345 68.935 77.515 69.105 ;
        RECT 77.805 68.935 77.975 69.105 ;
        RECT 78.265 68.935 78.435 69.105 ;
        RECT 78.725 68.935 78.895 69.105 ;
        RECT 79.185 68.935 79.355 69.105 ;
        RECT 79.645 68.935 79.815 69.105 ;
        RECT 80.105 68.935 80.275 69.105 ;
        RECT 80.565 68.935 80.735 69.105 ;
        RECT 81.025 68.935 81.195 69.105 ;
        RECT 81.485 68.935 81.655 69.105 ;
        RECT 81.945 68.935 82.115 69.105 ;
        RECT 82.405 68.935 82.575 69.105 ;
        RECT 82.865 68.935 83.035 69.105 ;
        RECT 83.325 68.935 83.495 69.105 ;
        RECT 83.785 68.935 83.955 69.105 ;
        RECT 84.245 68.935 84.415 69.105 ;
        RECT 84.705 68.935 84.875 69.105 ;
        RECT 85.165 68.935 85.335 69.105 ;
        RECT 85.625 68.935 85.795 69.105 ;
        RECT 86.085 68.935 86.255 69.105 ;
        RECT 86.545 68.935 86.715 69.105 ;
        RECT 87.005 68.935 87.175 69.105 ;
        RECT 87.465 68.935 87.635 69.105 ;
        RECT 87.925 68.935 88.095 69.105 ;
        RECT 88.385 68.935 88.555 69.105 ;
        RECT 88.845 68.935 89.015 69.105 ;
        RECT 89.305 68.935 89.475 69.105 ;
        RECT 89.765 68.935 89.935 69.105 ;
        RECT 90.225 68.935 90.395 69.105 ;
        RECT 90.685 68.935 90.855 69.105 ;
        RECT 91.145 68.935 91.315 69.105 ;
        RECT 91.605 68.935 91.775 69.105 ;
        RECT 92.065 68.935 92.235 69.105 ;
        RECT 92.525 68.935 92.695 69.105 ;
        RECT 92.985 68.935 93.155 69.105 ;
        RECT 93.445 68.935 93.615 69.105 ;
        RECT 93.905 68.935 94.075 69.105 ;
        RECT 94.365 68.935 94.535 69.105 ;
        RECT 94.825 68.935 94.995 69.105 ;
        RECT 95.285 68.935 95.455 69.105 ;
        RECT 95.745 68.935 95.915 69.105 ;
        RECT 96.205 68.935 96.375 69.105 ;
        RECT 96.665 68.935 96.835 69.105 ;
        RECT 97.125 68.935 97.295 69.105 ;
        RECT 97.585 68.935 97.755 69.105 ;
        RECT 98.045 68.935 98.215 69.105 ;
        RECT 98.505 68.935 98.675 69.105 ;
        RECT 98.965 68.935 99.135 69.105 ;
        RECT 99.425 68.935 99.595 69.105 ;
        RECT 99.885 68.935 100.055 69.105 ;
        RECT 100.345 68.935 100.515 69.105 ;
        RECT 100.805 68.935 100.975 69.105 ;
        RECT 101.265 68.935 101.435 69.105 ;
        RECT 101.725 68.935 101.895 69.105 ;
        RECT 102.185 68.935 102.355 69.105 ;
        RECT 102.645 68.935 102.815 69.105 ;
        RECT 103.105 68.935 103.275 69.105 ;
        RECT 103.565 68.935 103.735 69.105 ;
        RECT 104.025 68.935 104.195 69.105 ;
        RECT 104.485 68.935 104.655 69.105 ;
        RECT 104.945 68.935 105.115 69.105 ;
        RECT 105.405 68.935 105.575 69.105 ;
        RECT 105.865 68.935 106.035 69.105 ;
        RECT 106.325 68.935 106.495 69.105 ;
        RECT 106.785 68.935 106.955 69.105 ;
        RECT 107.245 68.935 107.415 69.105 ;
        RECT 107.705 68.935 107.875 69.105 ;
        RECT 108.165 68.935 108.335 69.105 ;
        RECT 108.625 68.935 108.795 69.105 ;
        RECT 109.085 68.935 109.255 69.105 ;
        RECT 109.545 68.935 109.715 69.105 ;
        RECT 110.005 68.935 110.175 69.105 ;
        RECT 110.465 68.935 110.635 69.105 ;
        RECT 110.925 68.935 111.095 69.105 ;
        RECT 111.385 68.935 111.555 69.105 ;
        RECT 111.845 68.935 112.015 69.105 ;
        RECT 112.305 68.935 112.475 69.105 ;
        RECT 112.765 68.935 112.935 69.105 ;
        RECT 113.225 68.935 113.395 69.105 ;
        RECT 113.685 68.935 113.855 69.105 ;
        RECT 114.145 68.935 114.315 69.105 ;
        RECT 114.605 68.935 114.775 69.105 ;
        RECT 115.065 68.935 115.235 69.105 ;
        RECT 115.525 68.935 115.695 69.105 ;
        RECT 115.985 68.935 116.155 69.105 ;
        RECT 116.445 68.935 116.615 69.105 ;
        RECT 116.905 68.935 117.075 69.105 ;
        RECT 117.365 68.935 117.535 69.105 ;
        RECT 117.825 68.935 117.995 69.105 ;
        RECT 118.285 68.935 118.455 69.105 ;
        RECT 118.745 68.935 118.915 69.105 ;
        RECT 119.205 68.935 119.375 69.105 ;
        RECT 119.665 68.935 119.835 69.105 ;
        RECT 120.125 68.935 120.295 69.105 ;
        RECT 120.585 68.935 120.755 69.105 ;
        RECT 121.045 68.935 121.215 69.105 ;
        RECT 121.505 68.935 121.675 69.105 ;
        RECT 121.965 68.935 122.135 69.105 ;
        RECT 122.425 68.935 122.595 69.105 ;
        RECT 122.885 68.935 123.055 69.105 ;
        RECT 123.345 68.935 123.515 69.105 ;
        RECT 123.805 68.935 123.975 69.105 ;
        RECT 124.265 68.935 124.435 69.105 ;
        RECT 124.725 68.935 124.895 69.105 ;
        RECT 125.185 68.935 125.355 69.105 ;
        RECT 125.645 68.935 125.815 69.105 ;
        RECT 126.105 68.935 126.275 69.105 ;
        RECT 126.565 68.935 126.735 69.105 ;
        RECT 127.025 68.935 127.195 69.105 ;
        RECT 127.485 68.935 127.655 69.105 ;
        RECT 127.945 68.935 128.115 69.105 ;
        RECT 128.405 68.935 128.575 69.105 ;
        RECT 128.865 68.935 129.035 69.105 ;
        RECT 129.325 68.935 129.495 69.105 ;
        RECT 129.785 68.935 129.955 69.105 ;
        RECT 130.245 68.935 130.415 69.105 ;
        RECT 130.705 68.935 130.875 69.105 ;
        RECT 131.165 68.935 131.335 69.105 ;
        RECT 131.625 68.935 131.795 69.105 ;
        RECT 132.085 68.935 132.255 69.105 ;
        RECT 132.545 68.935 132.715 69.105 ;
        RECT 133.005 68.935 133.175 69.105 ;
        RECT 133.465 68.935 133.635 69.105 ;
        RECT 133.925 68.935 134.095 69.105 ;
        RECT 134.385 68.935 134.555 69.105 ;
        RECT 134.845 68.935 135.015 69.105 ;
        RECT 135.305 68.935 135.475 69.105 ;
        RECT 135.765 68.935 135.935 69.105 ;
        RECT 136.225 68.935 136.395 69.105 ;
        RECT 136.685 68.935 136.855 69.105 ;
        RECT 137.145 68.935 137.315 69.105 ;
        RECT 137.605 68.935 137.775 69.105 ;
        RECT 138.065 68.935 138.235 69.105 ;
        RECT 138.525 68.935 138.695 69.105 ;
        RECT 138.985 68.935 139.155 69.105 ;
        RECT 50.665 66.215 50.835 66.385 ;
        RECT 51.125 66.215 51.295 66.385 ;
        RECT 51.585 66.215 51.755 66.385 ;
        RECT 52.045 66.215 52.215 66.385 ;
        RECT 52.505 66.215 52.675 66.385 ;
        RECT 52.965 66.215 53.135 66.385 ;
        RECT 53.425 66.215 53.595 66.385 ;
        RECT 53.885 66.215 54.055 66.385 ;
        RECT 54.345 66.215 54.515 66.385 ;
        RECT 54.805 66.215 54.975 66.385 ;
        RECT 55.265 66.215 55.435 66.385 ;
        RECT 55.725 66.215 55.895 66.385 ;
        RECT 56.185 66.215 56.355 66.385 ;
        RECT 56.645 66.215 56.815 66.385 ;
        RECT 57.105 66.215 57.275 66.385 ;
        RECT 57.565 66.215 57.735 66.385 ;
        RECT 58.025 66.215 58.195 66.385 ;
        RECT 58.485 66.215 58.655 66.385 ;
        RECT 58.945 66.215 59.115 66.385 ;
        RECT 59.405 66.215 59.575 66.385 ;
        RECT 59.865 66.215 60.035 66.385 ;
        RECT 60.325 66.215 60.495 66.385 ;
        RECT 60.785 66.215 60.955 66.385 ;
        RECT 61.245 66.215 61.415 66.385 ;
        RECT 61.705 66.215 61.875 66.385 ;
        RECT 62.165 66.215 62.335 66.385 ;
        RECT 62.625 66.215 62.795 66.385 ;
        RECT 63.085 66.215 63.255 66.385 ;
        RECT 63.545 66.215 63.715 66.385 ;
        RECT 64.005 66.215 64.175 66.385 ;
        RECT 64.465 66.215 64.635 66.385 ;
        RECT 64.925 66.215 65.095 66.385 ;
        RECT 65.385 66.215 65.555 66.385 ;
        RECT 65.845 66.215 66.015 66.385 ;
        RECT 66.305 66.215 66.475 66.385 ;
        RECT 66.765 66.215 66.935 66.385 ;
        RECT 67.225 66.215 67.395 66.385 ;
        RECT 67.685 66.215 67.855 66.385 ;
        RECT 68.145 66.215 68.315 66.385 ;
        RECT 68.605 66.215 68.775 66.385 ;
        RECT 69.065 66.215 69.235 66.385 ;
        RECT 69.525 66.215 69.695 66.385 ;
        RECT 69.985 66.215 70.155 66.385 ;
        RECT 70.445 66.215 70.615 66.385 ;
        RECT 70.905 66.215 71.075 66.385 ;
        RECT 71.365 66.215 71.535 66.385 ;
        RECT 71.825 66.215 71.995 66.385 ;
        RECT 72.285 66.215 72.455 66.385 ;
        RECT 72.745 66.215 72.915 66.385 ;
        RECT 73.205 66.215 73.375 66.385 ;
        RECT 73.665 66.215 73.835 66.385 ;
        RECT 74.125 66.215 74.295 66.385 ;
        RECT 74.585 66.215 74.755 66.385 ;
        RECT 75.045 66.215 75.215 66.385 ;
        RECT 75.505 66.215 75.675 66.385 ;
        RECT 75.965 66.215 76.135 66.385 ;
        RECT 76.425 66.215 76.595 66.385 ;
        RECT 76.885 66.215 77.055 66.385 ;
        RECT 77.345 66.215 77.515 66.385 ;
        RECT 77.805 66.215 77.975 66.385 ;
        RECT 78.265 66.215 78.435 66.385 ;
        RECT 78.725 66.215 78.895 66.385 ;
        RECT 79.185 66.215 79.355 66.385 ;
        RECT 79.645 66.215 79.815 66.385 ;
        RECT 80.105 66.215 80.275 66.385 ;
        RECT 80.565 66.215 80.735 66.385 ;
        RECT 81.025 66.215 81.195 66.385 ;
        RECT 81.485 66.215 81.655 66.385 ;
        RECT 81.945 66.215 82.115 66.385 ;
        RECT 82.405 66.215 82.575 66.385 ;
        RECT 82.865 66.215 83.035 66.385 ;
        RECT 83.325 66.215 83.495 66.385 ;
        RECT 83.785 66.215 83.955 66.385 ;
        RECT 84.245 66.215 84.415 66.385 ;
        RECT 84.705 66.215 84.875 66.385 ;
        RECT 85.165 66.215 85.335 66.385 ;
        RECT 85.625 66.215 85.795 66.385 ;
        RECT 86.085 66.215 86.255 66.385 ;
        RECT 86.545 66.215 86.715 66.385 ;
        RECT 87.005 66.215 87.175 66.385 ;
        RECT 87.465 66.215 87.635 66.385 ;
        RECT 87.925 66.215 88.095 66.385 ;
        RECT 88.385 66.215 88.555 66.385 ;
        RECT 88.845 66.215 89.015 66.385 ;
        RECT 89.305 66.215 89.475 66.385 ;
        RECT 89.765 66.215 89.935 66.385 ;
        RECT 90.225 66.215 90.395 66.385 ;
        RECT 90.685 66.215 90.855 66.385 ;
        RECT 91.145 66.215 91.315 66.385 ;
        RECT 91.605 66.215 91.775 66.385 ;
        RECT 92.065 66.215 92.235 66.385 ;
        RECT 92.525 66.215 92.695 66.385 ;
        RECT 92.985 66.215 93.155 66.385 ;
        RECT 93.445 66.215 93.615 66.385 ;
        RECT 93.905 66.215 94.075 66.385 ;
        RECT 94.365 66.215 94.535 66.385 ;
        RECT 94.825 66.215 94.995 66.385 ;
        RECT 95.285 66.215 95.455 66.385 ;
        RECT 95.745 66.215 95.915 66.385 ;
        RECT 96.205 66.215 96.375 66.385 ;
        RECT 96.665 66.215 96.835 66.385 ;
        RECT 97.125 66.215 97.295 66.385 ;
        RECT 97.585 66.215 97.755 66.385 ;
        RECT 98.045 66.215 98.215 66.385 ;
        RECT 98.505 66.215 98.675 66.385 ;
        RECT 98.965 66.215 99.135 66.385 ;
        RECT 99.425 66.215 99.595 66.385 ;
        RECT 99.885 66.215 100.055 66.385 ;
        RECT 100.345 66.215 100.515 66.385 ;
        RECT 100.805 66.215 100.975 66.385 ;
        RECT 101.265 66.215 101.435 66.385 ;
        RECT 101.725 66.215 101.895 66.385 ;
        RECT 102.185 66.215 102.355 66.385 ;
        RECT 102.645 66.215 102.815 66.385 ;
        RECT 103.105 66.215 103.275 66.385 ;
        RECT 103.565 66.215 103.735 66.385 ;
        RECT 104.025 66.215 104.195 66.385 ;
        RECT 104.485 66.215 104.655 66.385 ;
        RECT 104.945 66.215 105.115 66.385 ;
        RECT 105.405 66.215 105.575 66.385 ;
        RECT 105.865 66.215 106.035 66.385 ;
        RECT 106.325 66.215 106.495 66.385 ;
        RECT 106.785 66.215 106.955 66.385 ;
        RECT 107.245 66.215 107.415 66.385 ;
        RECT 107.705 66.215 107.875 66.385 ;
        RECT 108.165 66.215 108.335 66.385 ;
        RECT 108.625 66.215 108.795 66.385 ;
        RECT 109.085 66.215 109.255 66.385 ;
        RECT 109.545 66.215 109.715 66.385 ;
        RECT 110.005 66.215 110.175 66.385 ;
        RECT 110.465 66.215 110.635 66.385 ;
        RECT 110.925 66.215 111.095 66.385 ;
        RECT 111.385 66.215 111.555 66.385 ;
        RECT 111.845 66.215 112.015 66.385 ;
        RECT 112.305 66.215 112.475 66.385 ;
        RECT 112.765 66.215 112.935 66.385 ;
        RECT 113.225 66.215 113.395 66.385 ;
        RECT 113.685 66.215 113.855 66.385 ;
        RECT 114.145 66.215 114.315 66.385 ;
        RECT 114.605 66.215 114.775 66.385 ;
        RECT 115.065 66.215 115.235 66.385 ;
        RECT 115.525 66.215 115.695 66.385 ;
        RECT 115.985 66.215 116.155 66.385 ;
        RECT 116.445 66.215 116.615 66.385 ;
        RECT 116.905 66.215 117.075 66.385 ;
        RECT 117.365 66.215 117.535 66.385 ;
        RECT 117.825 66.215 117.995 66.385 ;
        RECT 118.285 66.215 118.455 66.385 ;
        RECT 118.745 66.215 118.915 66.385 ;
        RECT 119.205 66.215 119.375 66.385 ;
        RECT 119.665 66.215 119.835 66.385 ;
        RECT 120.125 66.215 120.295 66.385 ;
        RECT 120.585 66.215 120.755 66.385 ;
        RECT 121.045 66.215 121.215 66.385 ;
        RECT 121.505 66.215 121.675 66.385 ;
        RECT 121.965 66.215 122.135 66.385 ;
        RECT 122.425 66.215 122.595 66.385 ;
        RECT 122.885 66.215 123.055 66.385 ;
        RECT 123.345 66.215 123.515 66.385 ;
        RECT 123.805 66.215 123.975 66.385 ;
        RECT 124.265 66.215 124.435 66.385 ;
        RECT 124.725 66.215 124.895 66.385 ;
        RECT 125.185 66.215 125.355 66.385 ;
        RECT 125.645 66.215 125.815 66.385 ;
        RECT 126.105 66.215 126.275 66.385 ;
        RECT 126.565 66.215 126.735 66.385 ;
        RECT 127.025 66.215 127.195 66.385 ;
        RECT 127.485 66.215 127.655 66.385 ;
        RECT 127.945 66.215 128.115 66.385 ;
        RECT 128.405 66.215 128.575 66.385 ;
        RECT 128.865 66.215 129.035 66.385 ;
        RECT 129.325 66.215 129.495 66.385 ;
        RECT 129.785 66.215 129.955 66.385 ;
        RECT 130.245 66.215 130.415 66.385 ;
        RECT 130.705 66.215 130.875 66.385 ;
        RECT 131.165 66.215 131.335 66.385 ;
        RECT 131.625 66.215 131.795 66.385 ;
        RECT 132.085 66.215 132.255 66.385 ;
        RECT 132.545 66.215 132.715 66.385 ;
        RECT 133.005 66.215 133.175 66.385 ;
        RECT 133.465 66.215 133.635 66.385 ;
        RECT 133.925 66.215 134.095 66.385 ;
        RECT 134.385 66.215 134.555 66.385 ;
        RECT 134.845 66.215 135.015 66.385 ;
        RECT 135.305 66.215 135.475 66.385 ;
        RECT 135.765 66.215 135.935 66.385 ;
        RECT 136.225 66.215 136.395 66.385 ;
        RECT 136.685 66.215 136.855 66.385 ;
        RECT 137.145 66.215 137.315 66.385 ;
        RECT 137.605 66.215 137.775 66.385 ;
        RECT 138.065 66.215 138.235 66.385 ;
        RECT 138.525 66.215 138.695 66.385 ;
        RECT 138.985 66.215 139.155 66.385 ;
        RECT 50.665 63.495 50.835 63.665 ;
        RECT 51.125 63.495 51.295 63.665 ;
        RECT 51.585 63.495 51.755 63.665 ;
        RECT 52.045 63.495 52.215 63.665 ;
        RECT 52.505 63.495 52.675 63.665 ;
        RECT 52.965 63.495 53.135 63.665 ;
        RECT 53.425 63.495 53.595 63.665 ;
        RECT 53.885 63.495 54.055 63.665 ;
        RECT 54.345 63.495 54.515 63.665 ;
        RECT 54.805 63.495 54.975 63.665 ;
        RECT 55.265 63.495 55.435 63.665 ;
        RECT 55.725 63.495 55.895 63.665 ;
        RECT 56.185 63.495 56.355 63.665 ;
        RECT 56.645 63.495 56.815 63.665 ;
        RECT 57.105 63.495 57.275 63.665 ;
        RECT 57.565 63.495 57.735 63.665 ;
        RECT 58.025 63.495 58.195 63.665 ;
        RECT 58.485 63.495 58.655 63.665 ;
        RECT 58.945 63.495 59.115 63.665 ;
        RECT 59.405 63.495 59.575 63.665 ;
        RECT 59.865 63.495 60.035 63.665 ;
        RECT 60.325 63.495 60.495 63.665 ;
        RECT 60.785 63.495 60.955 63.665 ;
        RECT 61.245 63.495 61.415 63.665 ;
        RECT 61.705 63.495 61.875 63.665 ;
        RECT 62.165 63.495 62.335 63.665 ;
        RECT 62.625 63.495 62.795 63.665 ;
        RECT 63.085 63.495 63.255 63.665 ;
        RECT 63.545 63.495 63.715 63.665 ;
        RECT 64.005 63.495 64.175 63.665 ;
        RECT 64.465 63.495 64.635 63.665 ;
        RECT 64.925 63.495 65.095 63.665 ;
        RECT 65.385 63.495 65.555 63.665 ;
        RECT 65.845 63.495 66.015 63.665 ;
        RECT 66.305 63.495 66.475 63.665 ;
        RECT 66.765 63.495 66.935 63.665 ;
        RECT 67.225 63.495 67.395 63.665 ;
        RECT 67.685 63.495 67.855 63.665 ;
        RECT 68.145 63.495 68.315 63.665 ;
        RECT 68.605 63.495 68.775 63.665 ;
        RECT 69.065 63.495 69.235 63.665 ;
        RECT 69.525 63.495 69.695 63.665 ;
        RECT 69.985 63.495 70.155 63.665 ;
        RECT 70.445 63.495 70.615 63.665 ;
        RECT 70.905 63.495 71.075 63.665 ;
        RECT 71.365 63.495 71.535 63.665 ;
        RECT 71.825 63.495 71.995 63.665 ;
        RECT 72.285 63.495 72.455 63.665 ;
        RECT 72.745 63.495 72.915 63.665 ;
        RECT 73.205 63.495 73.375 63.665 ;
        RECT 73.665 63.495 73.835 63.665 ;
        RECT 74.125 63.495 74.295 63.665 ;
        RECT 74.585 63.495 74.755 63.665 ;
        RECT 75.045 63.495 75.215 63.665 ;
        RECT 75.505 63.495 75.675 63.665 ;
        RECT 75.965 63.495 76.135 63.665 ;
        RECT 76.425 63.495 76.595 63.665 ;
        RECT 76.885 63.495 77.055 63.665 ;
        RECT 77.345 63.495 77.515 63.665 ;
        RECT 77.805 63.495 77.975 63.665 ;
        RECT 78.265 63.495 78.435 63.665 ;
        RECT 78.725 63.495 78.895 63.665 ;
        RECT 79.185 63.495 79.355 63.665 ;
        RECT 79.645 63.495 79.815 63.665 ;
        RECT 80.105 63.495 80.275 63.665 ;
        RECT 80.565 63.495 80.735 63.665 ;
        RECT 81.025 63.495 81.195 63.665 ;
        RECT 81.485 63.495 81.655 63.665 ;
        RECT 81.945 63.495 82.115 63.665 ;
        RECT 82.405 63.495 82.575 63.665 ;
        RECT 82.865 63.495 83.035 63.665 ;
        RECT 83.325 63.495 83.495 63.665 ;
        RECT 83.785 63.495 83.955 63.665 ;
        RECT 84.245 63.495 84.415 63.665 ;
        RECT 84.705 63.495 84.875 63.665 ;
        RECT 85.165 63.495 85.335 63.665 ;
        RECT 85.625 63.495 85.795 63.665 ;
        RECT 86.085 63.495 86.255 63.665 ;
        RECT 86.545 63.495 86.715 63.665 ;
        RECT 87.005 63.495 87.175 63.665 ;
        RECT 87.465 63.495 87.635 63.665 ;
        RECT 87.925 63.495 88.095 63.665 ;
        RECT 88.385 63.495 88.555 63.665 ;
        RECT 88.845 63.495 89.015 63.665 ;
        RECT 89.305 63.495 89.475 63.665 ;
        RECT 89.765 63.495 89.935 63.665 ;
        RECT 90.225 63.495 90.395 63.665 ;
        RECT 90.685 63.495 90.855 63.665 ;
        RECT 91.145 63.495 91.315 63.665 ;
        RECT 91.605 63.495 91.775 63.665 ;
        RECT 92.065 63.495 92.235 63.665 ;
        RECT 92.525 63.495 92.695 63.665 ;
        RECT 92.985 63.495 93.155 63.665 ;
        RECT 93.445 63.495 93.615 63.665 ;
        RECT 93.905 63.495 94.075 63.665 ;
        RECT 94.365 63.495 94.535 63.665 ;
        RECT 94.825 63.495 94.995 63.665 ;
        RECT 95.285 63.495 95.455 63.665 ;
        RECT 95.745 63.495 95.915 63.665 ;
        RECT 96.205 63.495 96.375 63.665 ;
        RECT 96.665 63.495 96.835 63.665 ;
        RECT 97.125 63.495 97.295 63.665 ;
        RECT 97.585 63.495 97.755 63.665 ;
        RECT 98.045 63.495 98.215 63.665 ;
        RECT 98.505 63.495 98.675 63.665 ;
        RECT 98.965 63.495 99.135 63.665 ;
        RECT 99.425 63.495 99.595 63.665 ;
        RECT 99.885 63.495 100.055 63.665 ;
        RECT 100.345 63.495 100.515 63.665 ;
        RECT 100.805 63.495 100.975 63.665 ;
        RECT 101.265 63.495 101.435 63.665 ;
        RECT 101.725 63.495 101.895 63.665 ;
        RECT 102.185 63.495 102.355 63.665 ;
        RECT 102.645 63.495 102.815 63.665 ;
        RECT 103.105 63.495 103.275 63.665 ;
        RECT 103.565 63.495 103.735 63.665 ;
        RECT 104.025 63.495 104.195 63.665 ;
        RECT 104.485 63.495 104.655 63.665 ;
        RECT 104.945 63.495 105.115 63.665 ;
        RECT 105.405 63.495 105.575 63.665 ;
        RECT 105.865 63.495 106.035 63.665 ;
        RECT 106.325 63.495 106.495 63.665 ;
        RECT 106.785 63.495 106.955 63.665 ;
        RECT 107.245 63.495 107.415 63.665 ;
        RECT 107.705 63.495 107.875 63.665 ;
        RECT 108.165 63.495 108.335 63.665 ;
        RECT 108.625 63.495 108.795 63.665 ;
        RECT 109.085 63.495 109.255 63.665 ;
        RECT 109.545 63.495 109.715 63.665 ;
        RECT 110.005 63.495 110.175 63.665 ;
        RECT 110.465 63.495 110.635 63.665 ;
        RECT 110.925 63.495 111.095 63.665 ;
        RECT 111.385 63.495 111.555 63.665 ;
        RECT 111.845 63.495 112.015 63.665 ;
        RECT 112.305 63.495 112.475 63.665 ;
        RECT 112.765 63.495 112.935 63.665 ;
        RECT 113.225 63.495 113.395 63.665 ;
        RECT 113.685 63.495 113.855 63.665 ;
        RECT 114.145 63.495 114.315 63.665 ;
        RECT 114.605 63.495 114.775 63.665 ;
        RECT 115.065 63.495 115.235 63.665 ;
        RECT 115.525 63.495 115.695 63.665 ;
        RECT 115.985 63.495 116.155 63.665 ;
        RECT 116.445 63.495 116.615 63.665 ;
        RECT 116.905 63.495 117.075 63.665 ;
        RECT 117.365 63.495 117.535 63.665 ;
        RECT 117.825 63.495 117.995 63.665 ;
        RECT 118.285 63.495 118.455 63.665 ;
        RECT 118.745 63.495 118.915 63.665 ;
        RECT 119.205 63.495 119.375 63.665 ;
        RECT 119.665 63.495 119.835 63.665 ;
        RECT 120.125 63.495 120.295 63.665 ;
        RECT 120.585 63.495 120.755 63.665 ;
        RECT 121.045 63.495 121.215 63.665 ;
        RECT 121.505 63.495 121.675 63.665 ;
        RECT 121.965 63.495 122.135 63.665 ;
        RECT 122.425 63.495 122.595 63.665 ;
        RECT 122.885 63.495 123.055 63.665 ;
        RECT 123.345 63.495 123.515 63.665 ;
        RECT 123.805 63.495 123.975 63.665 ;
        RECT 124.265 63.495 124.435 63.665 ;
        RECT 124.725 63.495 124.895 63.665 ;
        RECT 125.185 63.495 125.355 63.665 ;
        RECT 125.645 63.495 125.815 63.665 ;
        RECT 126.105 63.495 126.275 63.665 ;
        RECT 126.565 63.495 126.735 63.665 ;
        RECT 127.025 63.495 127.195 63.665 ;
        RECT 127.485 63.495 127.655 63.665 ;
        RECT 127.945 63.495 128.115 63.665 ;
        RECT 128.405 63.495 128.575 63.665 ;
        RECT 128.865 63.495 129.035 63.665 ;
        RECT 129.325 63.495 129.495 63.665 ;
        RECT 129.785 63.495 129.955 63.665 ;
        RECT 130.245 63.495 130.415 63.665 ;
        RECT 130.705 63.495 130.875 63.665 ;
        RECT 131.165 63.495 131.335 63.665 ;
        RECT 131.625 63.495 131.795 63.665 ;
        RECT 132.085 63.495 132.255 63.665 ;
        RECT 132.545 63.495 132.715 63.665 ;
        RECT 133.005 63.495 133.175 63.665 ;
        RECT 133.465 63.495 133.635 63.665 ;
        RECT 133.925 63.495 134.095 63.665 ;
        RECT 134.385 63.495 134.555 63.665 ;
        RECT 134.845 63.495 135.015 63.665 ;
        RECT 135.305 63.495 135.475 63.665 ;
        RECT 135.765 63.495 135.935 63.665 ;
        RECT 136.225 63.495 136.395 63.665 ;
        RECT 136.685 63.495 136.855 63.665 ;
        RECT 137.145 63.495 137.315 63.665 ;
        RECT 137.605 63.495 137.775 63.665 ;
        RECT 138.065 63.495 138.235 63.665 ;
        RECT 138.525 63.495 138.695 63.665 ;
        RECT 138.985 63.495 139.155 63.665 ;
        RECT 50.665 60.775 50.835 60.945 ;
        RECT 51.125 60.775 51.295 60.945 ;
        RECT 51.585 60.775 51.755 60.945 ;
        RECT 52.045 60.775 52.215 60.945 ;
        RECT 52.505 60.775 52.675 60.945 ;
        RECT 52.965 60.775 53.135 60.945 ;
        RECT 53.425 60.775 53.595 60.945 ;
        RECT 53.885 60.775 54.055 60.945 ;
        RECT 54.345 60.775 54.515 60.945 ;
        RECT 54.805 60.775 54.975 60.945 ;
        RECT 55.265 60.775 55.435 60.945 ;
        RECT 55.725 60.775 55.895 60.945 ;
        RECT 56.185 60.775 56.355 60.945 ;
        RECT 56.645 60.775 56.815 60.945 ;
        RECT 57.105 60.775 57.275 60.945 ;
        RECT 57.565 60.775 57.735 60.945 ;
        RECT 58.025 60.775 58.195 60.945 ;
        RECT 58.485 60.775 58.655 60.945 ;
        RECT 58.945 60.775 59.115 60.945 ;
        RECT 59.405 60.775 59.575 60.945 ;
        RECT 59.865 60.775 60.035 60.945 ;
        RECT 60.325 60.775 60.495 60.945 ;
        RECT 60.785 60.775 60.955 60.945 ;
        RECT 61.245 60.775 61.415 60.945 ;
        RECT 61.705 60.775 61.875 60.945 ;
        RECT 62.165 60.775 62.335 60.945 ;
        RECT 62.625 60.775 62.795 60.945 ;
        RECT 63.085 60.775 63.255 60.945 ;
        RECT 63.545 60.775 63.715 60.945 ;
        RECT 64.005 60.775 64.175 60.945 ;
        RECT 64.465 60.775 64.635 60.945 ;
        RECT 64.925 60.775 65.095 60.945 ;
        RECT 65.385 60.775 65.555 60.945 ;
        RECT 65.845 60.775 66.015 60.945 ;
        RECT 66.305 60.775 66.475 60.945 ;
        RECT 66.765 60.775 66.935 60.945 ;
        RECT 67.225 60.775 67.395 60.945 ;
        RECT 67.685 60.775 67.855 60.945 ;
        RECT 68.145 60.775 68.315 60.945 ;
        RECT 68.605 60.775 68.775 60.945 ;
        RECT 69.065 60.775 69.235 60.945 ;
        RECT 69.525 60.775 69.695 60.945 ;
        RECT 69.985 60.775 70.155 60.945 ;
        RECT 70.445 60.775 70.615 60.945 ;
        RECT 70.905 60.775 71.075 60.945 ;
        RECT 71.365 60.775 71.535 60.945 ;
        RECT 71.825 60.775 71.995 60.945 ;
        RECT 72.285 60.775 72.455 60.945 ;
        RECT 72.745 60.775 72.915 60.945 ;
        RECT 73.205 60.775 73.375 60.945 ;
        RECT 73.665 60.775 73.835 60.945 ;
        RECT 74.125 60.775 74.295 60.945 ;
        RECT 74.585 60.775 74.755 60.945 ;
        RECT 75.045 60.775 75.215 60.945 ;
        RECT 75.505 60.775 75.675 60.945 ;
        RECT 75.965 60.775 76.135 60.945 ;
        RECT 76.425 60.775 76.595 60.945 ;
        RECT 76.885 60.775 77.055 60.945 ;
        RECT 77.345 60.775 77.515 60.945 ;
        RECT 77.805 60.775 77.975 60.945 ;
        RECT 78.265 60.775 78.435 60.945 ;
        RECT 78.725 60.775 78.895 60.945 ;
        RECT 79.185 60.775 79.355 60.945 ;
        RECT 79.645 60.775 79.815 60.945 ;
        RECT 80.105 60.775 80.275 60.945 ;
        RECT 80.565 60.775 80.735 60.945 ;
        RECT 81.025 60.775 81.195 60.945 ;
        RECT 81.485 60.775 81.655 60.945 ;
        RECT 81.945 60.775 82.115 60.945 ;
        RECT 82.405 60.775 82.575 60.945 ;
        RECT 82.865 60.775 83.035 60.945 ;
        RECT 83.325 60.775 83.495 60.945 ;
        RECT 83.785 60.775 83.955 60.945 ;
        RECT 84.245 60.775 84.415 60.945 ;
        RECT 84.705 60.775 84.875 60.945 ;
        RECT 85.165 60.775 85.335 60.945 ;
        RECT 85.625 60.775 85.795 60.945 ;
        RECT 86.085 60.775 86.255 60.945 ;
        RECT 86.545 60.775 86.715 60.945 ;
        RECT 87.005 60.775 87.175 60.945 ;
        RECT 87.465 60.775 87.635 60.945 ;
        RECT 87.925 60.775 88.095 60.945 ;
        RECT 88.385 60.775 88.555 60.945 ;
        RECT 88.845 60.775 89.015 60.945 ;
        RECT 89.305 60.775 89.475 60.945 ;
        RECT 89.765 60.775 89.935 60.945 ;
        RECT 90.225 60.775 90.395 60.945 ;
        RECT 90.685 60.775 90.855 60.945 ;
        RECT 91.145 60.775 91.315 60.945 ;
        RECT 91.605 60.775 91.775 60.945 ;
        RECT 92.065 60.775 92.235 60.945 ;
        RECT 92.525 60.775 92.695 60.945 ;
        RECT 92.985 60.775 93.155 60.945 ;
        RECT 93.445 60.775 93.615 60.945 ;
        RECT 93.905 60.775 94.075 60.945 ;
        RECT 94.365 60.775 94.535 60.945 ;
        RECT 94.825 60.775 94.995 60.945 ;
        RECT 95.285 60.775 95.455 60.945 ;
        RECT 95.745 60.775 95.915 60.945 ;
        RECT 96.205 60.775 96.375 60.945 ;
        RECT 96.665 60.775 96.835 60.945 ;
        RECT 97.125 60.775 97.295 60.945 ;
        RECT 97.585 60.775 97.755 60.945 ;
        RECT 98.045 60.775 98.215 60.945 ;
        RECT 98.505 60.775 98.675 60.945 ;
        RECT 98.965 60.775 99.135 60.945 ;
        RECT 99.425 60.775 99.595 60.945 ;
        RECT 99.885 60.775 100.055 60.945 ;
        RECT 100.345 60.775 100.515 60.945 ;
        RECT 100.805 60.775 100.975 60.945 ;
        RECT 101.265 60.775 101.435 60.945 ;
        RECT 101.725 60.775 101.895 60.945 ;
        RECT 102.185 60.775 102.355 60.945 ;
        RECT 102.645 60.775 102.815 60.945 ;
        RECT 103.105 60.775 103.275 60.945 ;
        RECT 103.565 60.775 103.735 60.945 ;
        RECT 104.025 60.775 104.195 60.945 ;
        RECT 104.485 60.775 104.655 60.945 ;
        RECT 104.945 60.775 105.115 60.945 ;
        RECT 105.405 60.775 105.575 60.945 ;
        RECT 105.865 60.775 106.035 60.945 ;
        RECT 106.325 60.775 106.495 60.945 ;
        RECT 106.785 60.775 106.955 60.945 ;
        RECT 107.245 60.775 107.415 60.945 ;
        RECT 107.705 60.775 107.875 60.945 ;
        RECT 108.165 60.775 108.335 60.945 ;
        RECT 108.625 60.775 108.795 60.945 ;
        RECT 109.085 60.775 109.255 60.945 ;
        RECT 109.545 60.775 109.715 60.945 ;
        RECT 110.005 60.775 110.175 60.945 ;
        RECT 110.465 60.775 110.635 60.945 ;
        RECT 110.925 60.775 111.095 60.945 ;
        RECT 111.385 60.775 111.555 60.945 ;
        RECT 111.845 60.775 112.015 60.945 ;
        RECT 112.305 60.775 112.475 60.945 ;
        RECT 112.765 60.775 112.935 60.945 ;
        RECT 113.225 60.775 113.395 60.945 ;
        RECT 113.685 60.775 113.855 60.945 ;
        RECT 114.145 60.775 114.315 60.945 ;
        RECT 114.605 60.775 114.775 60.945 ;
        RECT 115.065 60.775 115.235 60.945 ;
        RECT 115.525 60.775 115.695 60.945 ;
        RECT 115.985 60.775 116.155 60.945 ;
        RECT 116.445 60.775 116.615 60.945 ;
        RECT 116.905 60.775 117.075 60.945 ;
        RECT 117.365 60.775 117.535 60.945 ;
        RECT 117.825 60.775 117.995 60.945 ;
        RECT 118.285 60.775 118.455 60.945 ;
        RECT 118.745 60.775 118.915 60.945 ;
        RECT 119.205 60.775 119.375 60.945 ;
        RECT 119.665 60.775 119.835 60.945 ;
        RECT 120.125 60.775 120.295 60.945 ;
        RECT 120.585 60.775 120.755 60.945 ;
        RECT 121.045 60.775 121.215 60.945 ;
        RECT 121.505 60.775 121.675 60.945 ;
        RECT 121.965 60.775 122.135 60.945 ;
        RECT 122.425 60.775 122.595 60.945 ;
        RECT 122.885 60.775 123.055 60.945 ;
        RECT 123.345 60.775 123.515 60.945 ;
        RECT 123.805 60.775 123.975 60.945 ;
        RECT 124.265 60.775 124.435 60.945 ;
        RECT 124.725 60.775 124.895 60.945 ;
        RECT 125.185 60.775 125.355 60.945 ;
        RECT 125.645 60.775 125.815 60.945 ;
        RECT 126.105 60.775 126.275 60.945 ;
        RECT 126.565 60.775 126.735 60.945 ;
        RECT 127.025 60.775 127.195 60.945 ;
        RECT 127.485 60.775 127.655 60.945 ;
        RECT 127.945 60.775 128.115 60.945 ;
        RECT 128.405 60.775 128.575 60.945 ;
        RECT 128.865 60.775 129.035 60.945 ;
        RECT 129.325 60.775 129.495 60.945 ;
        RECT 129.785 60.775 129.955 60.945 ;
        RECT 130.245 60.775 130.415 60.945 ;
        RECT 130.705 60.775 130.875 60.945 ;
        RECT 131.165 60.775 131.335 60.945 ;
        RECT 131.625 60.775 131.795 60.945 ;
        RECT 132.085 60.775 132.255 60.945 ;
        RECT 132.545 60.775 132.715 60.945 ;
        RECT 133.005 60.775 133.175 60.945 ;
        RECT 133.465 60.775 133.635 60.945 ;
        RECT 133.925 60.775 134.095 60.945 ;
        RECT 134.385 60.775 134.555 60.945 ;
        RECT 134.845 60.775 135.015 60.945 ;
        RECT 135.305 60.775 135.475 60.945 ;
        RECT 135.765 60.775 135.935 60.945 ;
        RECT 136.225 60.775 136.395 60.945 ;
        RECT 136.685 60.775 136.855 60.945 ;
        RECT 137.145 60.775 137.315 60.945 ;
        RECT 137.605 60.775 137.775 60.945 ;
        RECT 138.065 60.775 138.235 60.945 ;
        RECT 138.525 60.775 138.695 60.945 ;
        RECT 138.985 60.775 139.155 60.945 ;
      LAYER met1 ;
        RECT 50.520 136.780 140.095 137.260 ;
        RECT 50.520 134.060 139.300 134.540 ;
        RECT 50.520 131.340 140.095 131.820 ;
        RECT 50.520 128.620 139.300 129.100 ;
        RECT 50.520 125.900 140.095 126.380 ;
        RECT 50.520 123.180 139.300 123.660 ;
        RECT 50.520 120.460 140.095 120.940 ;
        RECT 50.520 117.740 139.300 118.220 ;
        RECT 50.520 115.020 140.095 115.500 ;
        RECT 50.520 112.300 139.300 112.780 ;
        RECT 50.520 109.580 140.095 110.060 ;
        RECT 63.930 108.700 64.250 108.760 ;
        RECT 65.325 108.700 65.615 108.745 ;
        RECT 63.930 108.560 65.615 108.700 ;
        RECT 63.930 108.500 64.250 108.560 ;
        RECT 65.325 108.515 65.615 108.560 ;
        RECT 65.785 108.700 66.075 108.745 ;
        RECT 66.705 108.700 66.995 108.745 ;
        RECT 65.785 108.560 66.995 108.700 ;
        RECT 65.785 108.515 66.075 108.560 ;
        RECT 66.705 108.515 66.995 108.560 ;
        RECT 50.520 106.860 139.300 107.340 ;
        RECT 57.965 105.980 58.255 106.025 ;
        RECT 61.185 105.980 61.475 106.025 ;
        RECT 57.965 105.840 61.475 105.980 ;
        RECT 57.965 105.795 58.255 105.840 ;
        RECT 61.185 105.795 61.475 105.840 ;
        RECT 57.030 105.640 57.350 105.700 ;
        RECT 57.505 105.640 57.795 105.685 ;
        RECT 57.030 105.500 57.795 105.640 ;
        RECT 57.030 105.440 57.350 105.500 ;
        RECT 57.505 105.455 57.795 105.500 ;
        RECT 58.425 105.640 58.715 105.685 ;
        RECT 60.250 105.640 60.570 105.700 ;
        RECT 58.425 105.500 60.570 105.640 ;
        RECT 58.425 105.455 58.715 105.500 ;
        RECT 60.250 105.440 60.570 105.500 ;
        RECT 62.105 105.640 62.395 105.685 ;
        RECT 62.550 105.640 62.870 105.700 ;
        RECT 62.105 105.500 62.870 105.640 ;
        RECT 62.105 105.455 62.395 105.500 ;
        RECT 62.550 105.440 62.870 105.500 ;
        RECT 58.870 105.100 59.190 105.360 ;
        RECT 50.520 104.140 140.095 104.620 ;
        RECT 52.905 103.940 53.195 103.985 ;
        RECT 57.030 103.940 57.350 104.000 ;
        RECT 52.905 103.800 57.350 103.940 ;
        RECT 52.905 103.755 53.195 103.800 ;
        RECT 57.030 103.740 57.350 103.800 ;
        RECT 48.750 103.260 49.070 103.320 ;
        RECT 51.985 103.260 52.275 103.305 ;
        RECT 48.750 103.120 52.275 103.260 ;
        RECT 57.120 103.260 57.260 103.740 ;
        RECT 61.645 103.600 61.935 103.645 ;
        RECT 63.025 103.600 63.315 103.645 ;
        RECT 63.470 103.600 63.790 103.660 ;
        RECT 61.645 103.460 63.790 103.600 ;
        RECT 61.645 103.415 61.935 103.460 ;
        RECT 63.025 103.415 63.315 103.460 ;
        RECT 63.470 103.400 63.790 103.460 ;
        RECT 59.805 103.260 60.095 103.305 ;
        RECT 57.120 103.120 60.095 103.260 ;
        RECT 48.750 103.060 49.070 103.120 ;
        RECT 51.985 103.075 52.275 103.120 ;
        RECT 59.805 103.075 60.095 103.120 ;
        RECT 60.250 103.260 60.570 103.320 ;
        RECT 61.185 103.260 61.475 103.305 ;
        RECT 60.250 103.120 61.475 103.260 ;
        RECT 60.250 103.060 60.570 103.120 ;
        RECT 61.185 103.075 61.475 103.120 ;
        RECT 62.105 103.260 62.400 103.305 ;
        RECT 65.340 103.260 65.630 103.305 ;
        RECT 62.105 103.120 65.630 103.260 ;
        RECT 62.105 103.075 62.400 103.120 ;
        RECT 65.340 103.075 65.630 103.120 ;
        RECT 61.260 102.580 61.400 103.075 ;
        RECT 62.550 102.720 62.870 102.980 ;
        RECT 63.930 102.720 64.250 102.980 ;
        RECT 64.020 102.580 64.160 102.720 ;
        RECT 61.260 102.440 64.160 102.580 ;
        RECT 50.520 101.420 139.300 101.900 ;
        RECT 51.985 100.200 52.275 100.245 ;
        RECT 58.870 100.200 59.190 100.260 ;
        RECT 51.985 100.060 59.190 100.200 ;
        RECT 51.985 100.015 52.275 100.060 ;
        RECT 58.870 100.000 59.190 100.060 ;
        RECT 52.905 99.520 53.195 99.565 ;
        RECT 58.410 99.520 58.730 99.580 ;
        RECT 52.905 99.380 58.730 99.520 ;
        RECT 52.905 99.335 53.195 99.380 ;
        RECT 58.410 99.320 58.730 99.380 ;
        RECT 50.520 98.700 140.095 99.180 ;
        RECT 61.645 98.500 61.935 98.545 ;
        RECT 62.550 98.500 62.870 98.560 ;
        RECT 61.645 98.360 62.870 98.500 ;
        RECT 61.645 98.315 61.935 98.360 ;
        RECT 62.550 98.300 62.870 98.360 ;
        RECT 60.250 97.820 60.570 97.880 ;
        RECT 60.725 97.820 61.015 97.865 ;
        RECT 60.250 97.680 61.015 97.820 ;
        RECT 60.250 97.620 60.570 97.680 ;
        RECT 60.725 97.635 61.015 97.680 ;
        RECT 50.520 95.980 139.300 96.460 ;
        RECT 58.410 94.760 58.730 94.820 ;
        RECT 61.645 94.760 61.935 94.805 ;
        RECT 58.410 94.620 61.935 94.760 ;
        RECT 58.410 94.560 58.730 94.620 ;
        RECT 61.645 94.575 61.935 94.620 ;
        RECT 62.565 94.760 62.855 94.805 ;
        RECT 63.930 94.760 64.250 94.820 ;
        RECT 62.565 94.620 64.250 94.760 ;
        RECT 62.565 94.575 62.855 94.620 ;
        RECT 63.930 94.560 64.250 94.620 ;
        RECT 57.950 94.080 58.270 94.140 ;
        RECT 61.645 94.080 61.935 94.125 ;
        RECT 66.230 94.080 66.550 94.140 ;
        RECT 57.950 93.940 66.550 94.080 ;
        RECT 57.950 93.880 58.270 93.940 ;
        RECT 61.645 93.895 61.935 93.940 ;
        RECT 66.230 93.880 66.550 93.940 ;
        RECT 50.520 93.260 140.095 93.740 ;
        RECT 57.950 92.860 58.270 93.120 ;
        RECT 58.410 92.860 58.730 93.120 ;
        RECT 60.250 93.060 60.570 93.120 ;
        RECT 60.725 93.060 61.015 93.105 ;
        RECT 60.250 92.920 61.015 93.060 ;
        RECT 60.250 92.860 60.570 92.920 ;
        RECT 60.725 92.875 61.015 92.920 ;
        RECT 63.025 92.720 63.315 92.765 ;
        RECT 66.705 92.720 66.995 92.765 ;
        RECT 63.025 92.580 66.995 92.720 ;
        RECT 63.025 92.535 63.315 92.580 ;
        RECT 66.705 92.535 66.995 92.580 ;
        RECT 62.550 92.180 62.870 92.440 ;
        RECT 64.865 92.380 65.155 92.425 ;
        RECT 63.560 92.240 65.155 92.380 ;
        RECT 63.560 92.100 63.700 92.240 ;
        RECT 64.865 92.195 65.155 92.240 ;
        RECT 66.230 92.180 66.550 92.440 ;
        RECT 57.505 92.040 57.795 92.085 ;
        RECT 63.470 92.040 63.790 92.100 ;
        RECT 57.505 91.900 63.790 92.040 ;
        RECT 57.505 91.855 57.795 91.900 ;
        RECT 63.470 91.840 63.790 91.900 ;
        RECT 60.250 91.160 60.570 91.420 ;
        RECT 50.520 90.540 139.300 91.020 ;
        RECT 62.105 90.340 62.395 90.385 ;
        RECT 62.550 90.340 62.870 90.400 ;
        RECT 62.105 90.200 62.870 90.340 ;
        RECT 62.105 90.155 62.395 90.200 ;
        RECT 62.550 90.140 62.870 90.200 ;
        RECT 58.870 89.660 59.190 89.720 ;
        RECT 58.870 89.520 61.860 89.660 ;
        RECT 58.870 89.460 59.190 89.520 ;
        RECT 60.250 89.120 60.570 89.380 ;
        RECT 61.720 89.365 61.860 89.520 ;
        RECT 61.645 89.135 61.935 89.365 ;
        RECT 50.520 87.820 140.095 88.300 ;
        RECT 50.520 85.100 139.300 85.580 ;
        RECT 50.520 82.380 140.095 82.860 ;
        RECT 50.520 79.660 139.300 80.140 ;
        RECT 50.520 76.940 140.095 77.420 ;
        RECT 50.520 74.220 139.300 74.700 ;
        RECT 50.520 71.500 140.095 71.980 ;
        RECT 50.520 68.780 139.300 69.260 ;
        RECT 50.520 66.060 140.095 66.540 ;
        RECT 50.520 63.340 139.300 63.820 ;
        RECT 50.520 60.620 140.095 61.100 ;
      LAYER via ;
        RECT 71.940 136.890 72.200 137.150 ;
        RECT 72.260 136.890 72.520 137.150 ;
        RECT 72.580 136.890 72.840 137.150 ;
        RECT 72.900 136.890 73.160 137.150 ;
        RECT 73.220 136.890 73.480 137.150 ;
        RECT 94.135 136.890 94.395 137.150 ;
        RECT 94.455 136.890 94.715 137.150 ;
        RECT 94.775 136.890 95.035 137.150 ;
        RECT 95.095 136.890 95.355 137.150 ;
        RECT 95.415 136.890 95.675 137.150 ;
        RECT 116.330 136.890 116.590 137.150 ;
        RECT 116.650 136.890 116.910 137.150 ;
        RECT 116.970 136.890 117.230 137.150 ;
        RECT 117.290 136.890 117.550 137.150 ;
        RECT 117.610 136.890 117.870 137.150 ;
        RECT 138.525 136.890 138.785 137.150 ;
        RECT 138.845 136.890 139.105 137.150 ;
        RECT 139.165 136.890 139.425 137.150 ;
        RECT 139.485 136.890 139.745 137.150 ;
        RECT 139.805 136.890 140.065 137.150 ;
        RECT 60.845 134.170 61.105 134.430 ;
        RECT 61.165 134.170 61.425 134.430 ;
        RECT 61.485 134.170 61.745 134.430 ;
        RECT 61.805 134.170 62.065 134.430 ;
        RECT 62.125 134.170 62.385 134.430 ;
        RECT 83.040 134.170 83.300 134.430 ;
        RECT 83.360 134.170 83.620 134.430 ;
        RECT 83.680 134.170 83.940 134.430 ;
        RECT 84.000 134.170 84.260 134.430 ;
        RECT 84.320 134.170 84.580 134.430 ;
        RECT 105.235 134.170 105.495 134.430 ;
        RECT 105.555 134.170 105.815 134.430 ;
        RECT 105.875 134.170 106.135 134.430 ;
        RECT 106.195 134.170 106.455 134.430 ;
        RECT 106.515 134.170 106.775 134.430 ;
        RECT 127.430 134.170 127.690 134.430 ;
        RECT 127.750 134.170 128.010 134.430 ;
        RECT 128.070 134.170 128.330 134.430 ;
        RECT 128.390 134.170 128.650 134.430 ;
        RECT 128.710 134.170 128.970 134.430 ;
        RECT 71.940 131.450 72.200 131.710 ;
        RECT 72.260 131.450 72.520 131.710 ;
        RECT 72.580 131.450 72.840 131.710 ;
        RECT 72.900 131.450 73.160 131.710 ;
        RECT 73.220 131.450 73.480 131.710 ;
        RECT 94.135 131.450 94.395 131.710 ;
        RECT 94.455 131.450 94.715 131.710 ;
        RECT 94.775 131.450 95.035 131.710 ;
        RECT 95.095 131.450 95.355 131.710 ;
        RECT 95.415 131.450 95.675 131.710 ;
        RECT 116.330 131.450 116.590 131.710 ;
        RECT 116.650 131.450 116.910 131.710 ;
        RECT 116.970 131.450 117.230 131.710 ;
        RECT 117.290 131.450 117.550 131.710 ;
        RECT 117.610 131.450 117.870 131.710 ;
        RECT 138.525 131.450 138.785 131.710 ;
        RECT 138.845 131.450 139.105 131.710 ;
        RECT 139.165 131.450 139.425 131.710 ;
        RECT 139.485 131.450 139.745 131.710 ;
        RECT 139.805 131.450 140.065 131.710 ;
        RECT 60.845 128.730 61.105 128.990 ;
        RECT 61.165 128.730 61.425 128.990 ;
        RECT 61.485 128.730 61.745 128.990 ;
        RECT 61.805 128.730 62.065 128.990 ;
        RECT 62.125 128.730 62.385 128.990 ;
        RECT 83.040 128.730 83.300 128.990 ;
        RECT 83.360 128.730 83.620 128.990 ;
        RECT 83.680 128.730 83.940 128.990 ;
        RECT 84.000 128.730 84.260 128.990 ;
        RECT 84.320 128.730 84.580 128.990 ;
        RECT 105.235 128.730 105.495 128.990 ;
        RECT 105.555 128.730 105.815 128.990 ;
        RECT 105.875 128.730 106.135 128.990 ;
        RECT 106.195 128.730 106.455 128.990 ;
        RECT 106.515 128.730 106.775 128.990 ;
        RECT 127.430 128.730 127.690 128.990 ;
        RECT 127.750 128.730 128.010 128.990 ;
        RECT 128.070 128.730 128.330 128.990 ;
        RECT 128.390 128.730 128.650 128.990 ;
        RECT 128.710 128.730 128.970 128.990 ;
        RECT 71.940 126.010 72.200 126.270 ;
        RECT 72.260 126.010 72.520 126.270 ;
        RECT 72.580 126.010 72.840 126.270 ;
        RECT 72.900 126.010 73.160 126.270 ;
        RECT 73.220 126.010 73.480 126.270 ;
        RECT 94.135 126.010 94.395 126.270 ;
        RECT 94.455 126.010 94.715 126.270 ;
        RECT 94.775 126.010 95.035 126.270 ;
        RECT 95.095 126.010 95.355 126.270 ;
        RECT 95.415 126.010 95.675 126.270 ;
        RECT 116.330 126.010 116.590 126.270 ;
        RECT 116.650 126.010 116.910 126.270 ;
        RECT 116.970 126.010 117.230 126.270 ;
        RECT 117.290 126.010 117.550 126.270 ;
        RECT 117.610 126.010 117.870 126.270 ;
        RECT 138.525 126.010 138.785 126.270 ;
        RECT 138.845 126.010 139.105 126.270 ;
        RECT 139.165 126.010 139.425 126.270 ;
        RECT 139.485 126.010 139.745 126.270 ;
        RECT 139.805 126.010 140.065 126.270 ;
        RECT 60.845 123.290 61.105 123.550 ;
        RECT 61.165 123.290 61.425 123.550 ;
        RECT 61.485 123.290 61.745 123.550 ;
        RECT 61.805 123.290 62.065 123.550 ;
        RECT 62.125 123.290 62.385 123.550 ;
        RECT 83.040 123.290 83.300 123.550 ;
        RECT 83.360 123.290 83.620 123.550 ;
        RECT 83.680 123.290 83.940 123.550 ;
        RECT 84.000 123.290 84.260 123.550 ;
        RECT 84.320 123.290 84.580 123.550 ;
        RECT 105.235 123.290 105.495 123.550 ;
        RECT 105.555 123.290 105.815 123.550 ;
        RECT 105.875 123.290 106.135 123.550 ;
        RECT 106.195 123.290 106.455 123.550 ;
        RECT 106.515 123.290 106.775 123.550 ;
        RECT 127.430 123.290 127.690 123.550 ;
        RECT 127.750 123.290 128.010 123.550 ;
        RECT 128.070 123.290 128.330 123.550 ;
        RECT 128.390 123.290 128.650 123.550 ;
        RECT 128.710 123.290 128.970 123.550 ;
        RECT 71.940 120.570 72.200 120.830 ;
        RECT 72.260 120.570 72.520 120.830 ;
        RECT 72.580 120.570 72.840 120.830 ;
        RECT 72.900 120.570 73.160 120.830 ;
        RECT 73.220 120.570 73.480 120.830 ;
        RECT 94.135 120.570 94.395 120.830 ;
        RECT 94.455 120.570 94.715 120.830 ;
        RECT 94.775 120.570 95.035 120.830 ;
        RECT 95.095 120.570 95.355 120.830 ;
        RECT 95.415 120.570 95.675 120.830 ;
        RECT 116.330 120.570 116.590 120.830 ;
        RECT 116.650 120.570 116.910 120.830 ;
        RECT 116.970 120.570 117.230 120.830 ;
        RECT 117.290 120.570 117.550 120.830 ;
        RECT 117.610 120.570 117.870 120.830 ;
        RECT 138.525 120.570 138.785 120.830 ;
        RECT 138.845 120.570 139.105 120.830 ;
        RECT 139.165 120.570 139.425 120.830 ;
        RECT 139.485 120.570 139.745 120.830 ;
        RECT 139.805 120.570 140.065 120.830 ;
        RECT 60.845 117.850 61.105 118.110 ;
        RECT 61.165 117.850 61.425 118.110 ;
        RECT 61.485 117.850 61.745 118.110 ;
        RECT 61.805 117.850 62.065 118.110 ;
        RECT 62.125 117.850 62.385 118.110 ;
        RECT 83.040 117.850 83.300 118.110 ;
        RECT 83.360 117.850 83.620 118.110 ;
        RECT 83.680 117.850 83.940 118.110 ;
        RECT 84.000 117.850 84.260 118.110 ;
        RECT 84.320 117.850 84.580 118.110 ;
        RECT 105.235 117.850 105.495 118.110 ;
        RECT 105.555 117.850 105.815 118.110 ;
        RECT 105.875 117.850 106.135 118.110 ;
        RECT 106.195 117.850 106.455 118.110 ;
        RECT 106.515 117.850 106.775 118.110 ;
        RECT 127.430 117.850 127.690 118.110 ;
        RECT 127.750 117.850 128.010 118.110 ;
        RECT 128.070 117.850 128.330 118.110 ;
        RECT 128.390 117.850 128.650 118.110 ;
        RECT 128.710 117.850 128.970 118.110 ;
        RECT 71.940 115.130 72.200 115.390 ;
        RECT 72.260 115.130 72.520 115.390 ;
        RECT 72.580 115.130 72.840 115.390 ;
        RECT 72.900 115.130 73.160 115.390 ;
        RECT 73.220 115.130 73.480 115.390 ;
        RECT 94.135 115.130 94.395 115.390 ;
        RECT 94.455 115.130 94.715 115.390 ;
        RECT 94.775 115.130 95.035 115.390 ;
        RECT 95.095 115.130 95.355 115.390 ;
        RECT 95.415 115.130 95.675 115.390 ;
        RECT 116.330 115.130 116.590 115.390 ;
        RECT 116.650 115.130 116.910 115.390 ;
        RECT 116.970 115.130 117.230 115.390 ;
        RECT 117.290 115.130 117.550 115.390 ;
        RECT 117.610 115.130 117.870 115.390 ;
        RECT 138.525 115.130 138.785 115.390 ;
        RECT 138.845 115.130 139.105 115.390 ;
        RECT 139.165 115.130 139.425 115.390 ;
        RECT 139.485 115.130 139.745 115.390 ;
        RECT 139.805 115.130 140.065 115.390 ;
        RECT 60.845 112.410 61.105 112.670 ;
        RECT 61.165 112.410 61.425 112.670 ;
        RECT 61.485 112.410 61.745 112.670 ;
        RECT 61.805 112.410 62.065 112.670 ;
        RECT 62.125 112.410 62.385 112.670 ;
        RECT 83.040 112.410 83.300 112.670 ;
        RECT 83.360 112.410 83.620 112.670 ;
        RECT 83.680 112.410 83.940 112.670 ;
        RECT 84.000 112.410 84.260 112.670 ;
        RECT 84.320 112.410 84.580 112.670 ;
        RECT 105.235 112.410 105.495 112.670 ;
        RECT 105.555 112.410 105.815 112.670 ;
        RECT 105.875 112.410 106.135 112.670 ;
        RECT 106.195 112.410 106.455 112.670 ;
        RECT 106.515 112.410 106.775 112.670 ;
        RECT 127.430 112.410 127.690 112.670 ;
        RECT 127.750 112.410 128.010 112.670 ;
        RECT 128.070 112.410 128.330 112.670 ;
        RECT 128.390 112.410 128.650 112.670 ;
        RECT 128.710 112.410 128.970 112.670 ;
        RECT 71.940 109.690 72.200 109.950 ;
        RECT 72.260 109.690 72.520 109.950 ;
        RECT 72.580 109.690 72.840 109.950 ;
        RECT 72.900 109.690 73.160 109.950 ;
        RECT 73.220 109.690 73.480 109.950 ;
        RECT 94.135 109.690 94.395 109.950 ;
        RECT 94.455 109.690 94.715 109.950 ;
        RECT 94.775 109.690 95.035 109.950 ;
        RECT 95.095 109.690 95.355 109.950 ;
        RECT 95.415 109.690 95.675 109.950 ;
        RECT 116.330 109.690 116.590 109.950 ;
        RECT 116.650 109.690 116.910 109.950 ;
        RECT 116.970 109.690 117.230 109.950 ;
        RECT 117.290 109.690 117.550 109.950 ;
        RECT 117.610 109.690 117.870 109.950 ;
        RECT 138.525 109.690 138.785 109.950 ;
        RECT 138.845 109.690 139.105 109.950 ;
        RECT 139.165 109.690 139.425 109.950 ;
        RECT 139.485 109.690 139.745 109.950 ;
        RECT 139.805 109.690 140.065 109.950 ;
        RECT 63.960 108.500 64.220 108.760 ;
        RECT 60.845 106.970 61.105 107.230 ;
        RECT 61.165 106.970 61.425 107.230 ;
        RECT 61.485 106.970 61.745 107.230 ;
        RECT 61.805 106.970 62.065 107.230 ;
        RECT 62.125 106.970 62.385 107.230 ;
        RECT 83.040 106.970 83.300 107.230 ;
        RECT 83.360 106.970 83.620 107.230 ;
        RECT 83.680 106.970 83.940 107.230 ;
        RECT 84.000 106.970 84.260 107.230 ;
        RECT 84.320 106.970 84.580 107.230 ;
        RECT 105.235 106.970 105.495 107.230 ;
        RECT 105.555 106.970 105.815 107.230 ;
        RECT 105.875 106.970 106.135 107.230 ;
        RECT 106.195 106.970 106.455 107.230 ;
        RECT 106.515 106.970 106.775 107.230 ;
        RECT 127.430 106.970 127.690 107.230 ;
        RECT 127.750 106.970 128.010 107.230 ;
        RECT 128.070 106.970 128.330 107.230 ;
        RECT 128.390 106.970 128.650 107.230 ;
        RECT 128.710 106.970 128.970 107.230 ;
        RECT 57.060 105.440 57.320 105.700 ;
        RECT 60.280 105.440 60.540 105.700 ;
        RECT 62.580 105.440 62.840 105.700 ;
        RECT 58.900 105.100 59.160 105.360 ;
        RECT 71.940 104.250 72.200 104.510 ;
        RECT 72.260 104.250 72.520 104.510 ;
        RECT 72.580 104.250 72.840 104.510 ;
        RECT 72.900 104.250 73.160 104.510 ;
        RECT 73.220 104.250 73.480 104.510 ;
        RECT 94.135 104.250 94.395 104.510 ;
        RECT 94.455 104.250 94.715 104.510 ;
        RECT 94.775 104.250 95.035 104.510 ;
        RECT 95.095 104.250 95.355 104.510 ;
        RECT 95.415 104.250 95.675 104.510 ;
        RECT 116.330 104.250 116.590 104.510 ;
        RECT 116.650 104.250 116.910 104.510 ;
        RECT 116.970 104.250 117.230 104.510 ;
        RECT 117.290 104.250 117.550 104.510 ;
        RECT 117.610 104.250 117.870 104.510 ;
        RECT 138.525 104.250 138.785 104.510 ;
        RECT 138.845 104.250 139.105 104.510 ;
        RECT 139.165 104.250 139.425 104.510 ;
        RECT 139.485 104.250 139.745 104.510 ;
        RECT 139.805 104.250 140.065 104.510 ;
        RECT 57.060 103.740 57.320 104.000 ;
        RECT 48.780 103.060 49.040 103.320 ;
        RECT 63.500 103.400 63.760 103.660 ;
        RECT 60.280 103.060 60.540 103.320 ;
        RECT 62.580 102.720 62.840 102.980 ;
        RECT 63.960 102.720 64.220 102.980 ;
        RECT 60.845 101.530 61.105 101.790 ;
        RECT 61.165 101.530 61.425 101.790 ;
        RECT 61.485 101.530 61.745 101.790 ;
        RECT 61.805 101.530 62.065 101.790 ;
        RECT 62.125 101.530 62.385 101.790 ;
        RECT 83.040 101.530 83.300 101.790 ;
        RECT 83.360 101.530 83.620 101.790 ;
        RECT 83.680 101.530 83.940 101.790 ;
        RECT 84.000 101.530 84.260 101.790 ;
        RECT 84.320 101.530 84.580 101.790 ;
        RECT 105.235 101.530 105.495 101.790 ;
        RECT 105.555 101.530 105.815 101.790 ;
        RECT 105.875 101.530 106.135 101.790 ;
        RECT 106.195 101.530 106.455 101.790 ;
        RECT 106.515 101.530 106.775 101.790 ;
        RECT 127.430 101.530 127.690 101.790 ;
        RECT 127.750 101.530 128.010 101.790 ;
        RECT 128.070 101.530 128.330 101.790 ;
        RECT 128.390 101.530 128.650 101.790 ;
        RECT 128.710 101.530 128.970 101.790 ;
        RECT 58.900 100.000 59.160 100.260 ;
        RECT 58.440 99.320 58.700 99.580 ;
        RECT 71.940 98.810 72.200 99.070 ;
        RECT 72.260 98.810 72.520 99.070 ;
        RECT 72.580 98.810 72.840 99.070 ;
        RECT 72.900 98.810 73.160 99.070 ;
        RECT 73.220 98.810 73.480 99.070 ;
        RECT 94.135 98.810 94.395 99.070 ;
        RECT 94.455 98.810 94.715 99.070 ;
        RECT 94.775 98.810 95.035 99.070 ;
        RECT 95.095 98.810 95.355 99.070 ;
        RECT 95.415 98.810 95.675 99.070 ;
        RECT 116.330 98.810 116.590 99.070 ;
        RECT 116.650 98.810 116.910 99.070 ;
        RECT 116.970 98.810 117.230 99.070 ;
        RECT 117.290 98.810 117.550 99.070 ;
        RECT 117.610 98.810 117.870 99.070 ;
        RECT 138.525 98.810 138.785 99.070 ;
        RECT 138.845 98.810 139.105 99.070 ;
        RECT 139.165 98.810 139.425 99.070 ;
        RECT 139.485 98.810 139.745 99.070 ;
        RECT 139.805 98.810 140.065 99.070 ;
        RECT 62.580 98.300 62.840 98.560 ;
        RECT 60.280 97.620 60.540 97.880 ;
        RECT 60.845 96.090 61.105 96.350 ;
        RECT 61.165 96.090 61.425 96.350 ;
        RECT 61.485 96.090 61.745 96.350 ;
        RECT 61.805 96.090 62.065 96.350 ;
        RECT 62.125 96.090 62.385 96.350 ;
        RECT 83.040 96.090 83.300 96.350 ;
        RECT 83.360 96.090 83.620 96.350 ;
        RECT 83.680 96.090 83.940 96.350 ;
        RECT 84.000 96.090 84.260 96.350 ;
        RECT 84.320 96.090 84.580 96.350 ;
        RECT 105.235 96.090 105.495 96.350 ;
        RECT 105.555 96.090 105.815 96.350 ;
        RECT 105.875 96.090 106.135 96.350 ;
        RECT 106.195 96.090 106.455 96.350 ;
        RECT 106.515 96.090 106.775 96.350 ;
        RECT 127.430 96.090 127.690 96.350 ;
        RECT 127.750 96.090 128.010 96.350 ;
        RECT 128.070 96.090 128.330 96.350 ;
        RECT 128.390 96.090 128.650 96.350 ;
        RECT 128.710 96.090 128.970 96.350 ;
        RECT 58.440 94.560 58.700 94.820 ;
        RECT 63.960 94.560 64.220 94.820 ;
        RECT 57.980 93.880 58.240 94.140 ;
        RECT 66.260 93.880 66.520 94.140 ;
        RECT 71.940 93.370 72.200 93.630 ;
        RECT 72.260 93.370 72.520 93.630 ;
        RECT 72.580 93.370 72.840 93.630 ;
        RECT 72.900 93.370 73.160 93.630 ;
        RECT 73.220 93.370 73.480 93.630 ;
        RECT 94.135 93.370 94.395 93.630 ;
        RECT 94.455 93.370 94.715 93.630 ;
        RECT 94.775 93.370 95.035 93.630 ;
        RECT 95.095 93.370 95.355 93.630 ;
        RECT 95.415 93.370 95.675 93.630 ;
        RECT 116.330 93.370 116.590 93.630 ;
        RECT 116.650 93.370 116.910 93.630 ;
        RECT 116.970 93.370 117.230 93.630 ;
        RECT 117.290 93.370 117.550 93.630 ;
        RECT 117.610 93.370 117.870 93.630 ;
        RECT 138.525 93.370 138.785 93.630 ;
        RECT 138.845 93.370 139.105 93.630 ;
        RECT 139.165 93.370 139.425 93.630 ;
        RECT 139.485 93.370 139.745 93.630 ;
        RECT 139.805 93.370 140.065 93.630 ;
        RECT 57.980 92.860 58.240 93.120 ;
        RECT 58.440 92.860 58.700 93.120 ;
        RECT 60.280 92.860 60.540 93.120 ;
        RECT 62.580 92.180 62.840 92.440 ;
        RECT 66.260 92.180 66.520 92.440 ;
        RECT 63.500 91.840 63.760 92.100 ;
        RECT 60.280 91.160 60.540 91.420 ;
        RECT 60.845 90.650 61.105 90.910 ;
        RECT 61.165 90.650 61.425 90.910 ;
        RECT 61.485 90.650 61.745 90.910 ;
        RECT 61.805 90.650 62.065 90.910 ;
        RECT 62.125 90.650 62.385 90.910 ;
        RECT 83.040 90.650 83.300 90.910 ;
        RECT 83.360 90.650 83.620 90.910 ;
        RECT 83.680 90.650 83.940 90.910 ;
        RECT 84.000 90.650 84.260 90.910 ;
        RECT 84.320 90.650 84.580 90.910 ;
        RECT 105.235 90.650 105.495 90.910 ;
        RECT 105.555 90.650 105.815 90.910 ;
        RECT 105.875 90.650 106.135 90.910 ;
        RECT 106.195 90.650 106.455 90.910 ;
        RECT 106.515 90.650 106.775 90.910 ;
        RECT 127.430 90.650 127.690 90.910 ;
        RECT 127.750 90.650 128.010 90.910 ;
        RECT 128.070 90.650 128.330 90.910 ;
        RECT 128.390 90.650 128.650 90.910 ;
        RECT 128.710 90.650 128.970 90.910 ;
        RECT 62.580 90.140 62.840 90.400 ;
        RECT 58.900 89.460 59.160 89.720 ;
        RECT 60.280 89.120 60.540 89.380 ;
        RECT 71.940 87.930 72.200 88.190 ;
        RECT 72.260 87.930 72.520 88.190 ;
        RECT 72.580 87.930 72.840 88.190 ;
        RECT 72.900 87.930 73.160 88.190 ;
        RECT 73.220 87.930 73.480 88.190 ;
        RECT 94.135 87.930 94.395 88.190 ;
        RECT 94.455 87.930 94.715 88.190 ;
        RECT 94.775 87.930 95.035 88.190 ;
        RECT 95.095 87.930 95.355 88.190 ;
        RECT 95.415 87.930 95.675 88.190 ;
        RECT 116.330 87.930 116.590 88.190 ;
        RECT 116.650 87.930 116.910 88.190 ;
        RECT 116.970 87.930 117.230 88.190 ;
        RECT 117.290 87.930 117.550 88.190 ;
        RECT 117.610 87.930 117.870 88.190 ;
        RECT 138.525 87.930 138.785 88.190 ;
        RECT 138.845 87.930 139.105 88.190 ;
        RECT 139.165 87.930 139.425 88.190 ;
        RECT 139.485 87.930 139.745 88.190 ;
        RECT 139.805 87.930 140.065 88.190 ;
        RECT 60.845 85.210 61.105 85.470 ;
        RECT 61.165 85.210 61.425 85.470 ;
        RECT 61.485 85.210 61.745 85.470 ;
        RECT 61.805 85.210 62.065 85.470 ;
        RECT 62.125 85.210 62.385 85.470 ;
        RECT 83.040 85.210 83.300 85.470 ;
        RECT 83.360 85.210 83.620 85.470 ;
        RECT 83.680 85.210 83.940 85.470 ;
        RECT 84.000 85.210 84.260 85.470 ;
        RECT 84.320 85.210 84.580 85.470 ;
        RECT 105.235 85.210 105.495 85.470 ;
        RECT 105.555 85.210 105.815 85.470 ;
        RECT 105.875 85.210 106.135 85.470 ;
        RECT 106.195 85.210 106.455 85.470 ;
        RECT 106.515 85.210 106.775 85.470 ;
        RECT 127.430 85.210 127.690 85.470 ;
        RECT 127.750 85.210 128.010 85.470 ;
        RECT 128.070 85.210 128.330 85.470 ;
        RECT 128.390 85.210 128.650 85.470 ;
        RECT 128.710 85.210 128.970 85.470 ;
        RECT 71.940 82.490 72.200 82.750 ;
        RECT 72.260 82.490 72.520 82.750 ;
        RECT 72.580 82.490 72.840 82.750 ;
        RECT 72.900 82.490 73.160 82.750 ;
        RECT 73.220 82.490 73.480 82.750 ;
        RECT 94.135 82.490 94.395 82.750 ;
        RECT 94.455 82.490 94.715 82.750 ;
        RECT 94.775 82.490 95.035 82.750 ;
        RECT 95.095 82.490 95.355 82.750 ;
        RECT 95.415 82.490 95.675 82.750 ;
        RECT 116.330 82.490 116.590 82.750 ;
        RECT 116.650 82.490 116.910 82.750 ;
        RECT 116.970 82.490 117.230 82.750 ;
        RECT 117.290 82.490 117.550 82.750 ;
        RECT 117.610 82.490 117.870 82.750 ;
        RECT 138.525 82.490 138.785 82.750 ;
        RECT 138.845 82.490 139.105 82.750 ;
        RECT 139.165 82.490 139.425 82.750 ;
        RECT 139.485 82.490 139.745 82.750 ;
        RECT 139.805 82.490 140.065 82.750 ;
        RECT 60.845 79.770 61.105 80.030 ;
        RECT 61.165 79.770 61.425 80.030 ;
        RECT 61.485 79.770 61.745 80.030 ;
        RECT 61.805 79.770 62.065 80.030 ;
        RECT 62.125 79.770 62.385 80.030 ;
        RECT 83.040 79.770 83.300 80.030 ;
        RECT 83.360 79.770 83.620 80.030 ;
        RECT 83.680 79.770 83.940 80.030 ;
        RECT 84.000 79.770 84.260 80.030 ;
        RECT 84.320 79.770 84.580 80.030 ;
        RECT 105.235 79.770 105.495 80.030 ;
        RECT 105.555 79.770 105.815 80.030 ;
        RECT 105.875 79.770 106.135 80.030 ;
        RECT 106.195 79.770 106.455 80.030 ;
        RECT 106.515 79.770 106.775 80.030 ;
        RECT 127.430 79.770 127.690 80.030 ;
        RECT 127.750 79.770 128.010 80.030 ;
        RECT 128.070 79.770 128.330 80.030 ;
        RECT 128.390 79.770 128.650 80.030 ;
        RECT 128.710 79.770 128.970 80.030 ;
        RECT 71.940 77.050 72.200 77.310 ;
        RECT 72.260 77.050 72.520 77.310 ;
        RECT 72.580 77.050 72.840 77.310 ;
        RECT 72.900 77.050 73.160 77.310 ;
        RECT 73.220 77.050 73.480 77.310 ;
        RECT 94.135 77.050 94.395 77.310 ;
        RECT 94.455 77.050 94.715 77.310 ;
        RECT 94.775 77.050 95.035 77.310 ;
        RECT 95.095 77.050 95.355 77.310 ;
        RECT 95.415 77.050 95.675 77.310 ;
        RECT 116.330 77.050 116.590 77.310 ;
        RECT 116.650 77.050 116.910 77.310 ;
        RECT 116.970 77.050 117.230 77.310 ;
        RECT 117.290 77.050 117.550 77.310 ;
        RECT 117.610 77.050 117.870 77.310 ;
        RECT 138.525 77.050 138.785 77.310 ;
        RECT 138.845 77.050 139.105 77.310 ;
        RECT 139.165 77.050 139.425 77.310 ;
        RECT 139.485 77.050 139.745 77.310 ;
        RECT 139.805 77.050 140.065 77.310 ;
        RECT 60.845 74.330 61.105 74.590 ;
        RECT 61.165 74.330 61.425 74.590 ;
        RECT 61.485 74.330 61.745 74.590 ;
        RECT 61.805 74.330 62.065 74.590 ;
        RECT 62.125 74.330 62.385 74.590 ;
        RECT 83.040 74.330 83.300 74.590 ;
        RECT 83.360 74.330 83.620 74.590 ;
        RECT 83.680 74.330 83.940 74.590 ;
        RECT 84.000 74.330 84.260 74.590 ;
        RECT 84.320 74.330 84.580 74.590 ;
        RECT 105.235 74.330 105.495 74.590 ;
        RECT 105.555 74.330 105.815 74.590 ;
        RECT 105.875 74.330 106.135 74.590 ;
        RECT 106.195 74.330 106.455 74.590 ;
        RECT 106.515 74.330 106.775 74.590 ;
        RECT 127.430 74.330 127.690 74.590 ;
        RECT 127.750 74.330 128.010 74.590 ;
        RECT 128.070 74.330 128.330 74.590 ;
        RECT 128.390 74.330 128.650 74.590 ;
        RECT 128.710 74.330 128.970 74.590 ;
        RECT 71.940 71.610 72.200 71.870 ;
        RECT 72.260 71.610 72.520 71.870 ;
        RECT 72.580 71.610 72.840 71.870 ;
        RECT 72.900 71.610 73.160 71.870 ;
        RECT 73.220 71.610 73.480 71.870 ;
        RECT 94.135 71.610 94.395 71.870 ;
        RECT 94.455 71.610 94.715 71.870 ;
        RECT 94.775 71.610 95.035 71.870 ;
        RECT 95.095 71.610 95.355 71.870 ;
        RECT 95.415 71.610 95.675 71.870 ;
        RECT 116.330 71.610 116.590 71.870 ;
        RECT 116.650 71.610 116.910 71.870 ;
        RECT 116.970 71.610 117.230 71.870 ;
        RECT 117.290 71.610 117.550 71.870 ;
        RECT 117.610 71.610 117.870 71.870 ;
        RECT 138.525 71.610 138.785 71.870 ;
        RECT 138.845 71.610 139.105 71.870 ;
        RECT 139.165 71.610 139.425 71.870 ;
        RECT 139.485 71.610 139.745 71.870 ;
        RECT 139.805 71.610 140.065 71.870 ;
        RECT 60.845 68.890 61.105 69.150 ;
        RECT 61.165 68.890 61.425 69.150 ;
        RECT 61.485 68.890 61.745 69.150 ;
        RECT 61.805 68.890 62.065 69.150 ;
        RECT 62.125 68.890 62.385 69.150 ;
        RECT 83.040 68.890 83.300 69.150 ;
        RECT 83.360 68.890 83.620 69.150 ;
        RECT 83.680 68.890 83.940 69.150 ;
        RECT 84.000 68.890 84.260 69.150 ;
        RECT 84.320 68.890 84.580 69.150 ;
        RECT 105.235 68.890 105.495 69.150 ;
        RECT 105.555 68.890 105.815 69.150 ;
        RECT 105.875 68.890 106.135 69.150 ;
        RECT 106.195 68.890 106.455 69.150 ;
        RECT 106.515 68.890 106.775 69.150 ;
        RECT 127.430 68.890 127.690 69.150 ;
        RECT 127.750 68.890 128.010 69.150 ;
        RECT 128.070 68.890 128.330 69.150 ;
        RECT 128.390 68.890 128.650 69.150 ;
        RECT 128.710 68.890 128.970 69.150 ;
        RECT 71.940 66.170 72.200 66.430 ;
        RECT 72.260 66.170 72.520 66.430 ;
        RECT 72.580 66.170 72.840 66.430 ;
        RECT 72.900 66.170 73.160 66.430 ;
        RECT 73.220 66.170 73.480 66.430 ;
        RECT 94.135 66.170 94.395 66.430 ;
        RECT 94.455 66.170 94.715 66.430 ;
        RECT 94.775 66.170 95.035 66.430 ;
        RECT 95.095 66.170 95.355 66.430 ;
        RECT 95.415 66.170 95.675 66.430 ;
        RECT 116.330 66.170 116.590 66.430 ;
        RECT 116.650 66.170 116.910 66.430 ;
        RECT 116.970 66.170 117.230 66.430 ;
        RECT 117.290 66.170 117.550 66.430 ;
        RECT 117.610 66.170 117.870 66.430 ;
        RECT 138.525 66.170 138.785 66.430 ;
        RECT 138.845 66.170 139.105 66.430 ;
        RECT 139.165 66.170 139.425 66.430 ;
        RECT 139.485 66.170 139.745 66.430 ;
        RECT 139.805 66.170 140.065 66.430 ;
        RECT 60.845 63.450 61.105 63.710 ;
        RECT 61.165 63.450 61.425 63.710 ;
        RECT 61.485 63.450 61.745 63.710 ;
        RECT 61.805 63.450 62.065 63.710 ;
        RECT 62.125 63.450 62.385 63.710 ;
        RECT 83.040 63.450 83.300 63.710 ;
        RECT 83.360 63.450 83.620 63.710 ;
        RECT 83.680 63.450 83.940 63.710 ;
        RECT 84.000 63.450 84.260 63.710 ;
        RECT 84.320 63.450 84.580 63.710 ;
        RECT 105.235 63.450 105.495 63.710 ;
        RECT 105.555 63.450 105.815 63.710 ;
        RECT 105.875 63.450 106.135 63.710 ;
        RECT 106.195 63.450 106.455 63.710 ;
        RECT 106.515 63.450 106.775 63.710 ;
        RECT 127.430 63.450 127.690 63.710 ;
        RECT 127.750 63.450 128.010 63.710 ;
        RECT 128.070 63.450 128.330 63.710 ;
        RECT 128.390 63.450 128.650 63.710 ;
        RECT 128.710 63.450 128.970 63.710 ;
        RECT 71.940 60.730 72.200 60.990 ;
        RECT 72.260 60.730 72.520 60.990 ;
        RECT 72.580 60.730 72.840 60.990 ;
        RECT 72.900 60.730 73.160 60.990 ;
        RECT 73.220 60.730 73.480 60.990 ;
        RECT 94.135 60.730 94.395 60.990 ;
        RECT 94.455 60.730 94.715 60.990 ;
        RECT 94.775 60.730 95.035 60.990 ;
        RECT 95.095 60.730 95.355 60.990 ;
        RECT 95.415 60.730 95.675 60.990 ;
        RECT 116.330 60.730 116.590 60.990 ;
        RECT 116.650 60.730 116.910 60.990 ;
        RECT 116.970 60.730 117.230 60.990 ;
        RECT 117.290 60.730 117.550 60.990 ;
        RECT 117.610 60.730 117.870 60.990 ;
        RECT 138.525 60.730 138.785 60.990 ;
        RECT 138.845 60.730 139.105 60.990 ;
        RECT 139.165 60.730 139.425 60.990 ;
        RECT 139.485 60.730 139.745 60.990 ;
        RECT 139.805 60.730 140.065 60.990 ;
      LAYER met2 ;
        RECT 71.940 136.835 73.480 137.205 ;
        RECT 94.135 136.835 95.675 137.205 ;
        RECT 116.330 136.835 117.870 137.205 ;
        RECT 138.525 136.835 140.065 137.205 ;
        RECT 60.845 134.115 62.385 134.485 ;
        RECT 83.040 134.115 84.580 134.485 ;
        RECT 105.235 134.115 106.775 134.485 ;
        RECT 127.430 134.115 128.970 134.485 ;
        RECT 71.940 131.395 73.480 131.765 ;
        RECT 94.135 131.395 95.675 131.765 ;
        RECT 116.330 131.395 117.870 131.765 ;
        RECT 138.525 131.395 140.065 131.765 ;
        RECT 60.845 128.675 62.385 129.045 ;
        RECT 83.040 128.675 84.580 129.045 ;
        RECT 105.235 128.675 106.775 129.045 ;
        RECT 127.430 128.675 128.970 129.045 ;
        RECT 71.940 125.955 73.480 126.325 ;
        RECT 94.135 125.955 95.675 126.325 ;
        RECT 116.330 125.955 117.870 126.325 ;
        RECT 138.525 125.955 140.065 126.325 ;
        RECT 60.845 123.235 62.385 123.605 ;
        RECT 83.040 123.235 84.580 123.605 ;
        RECT 105.235 123.235 106.775 123.605 ;
        RECT 127.430 123.235 128.970 123.605 ;
        RECT 71.940 120.515 73.480 120.885 ;
        RECT 94.135 120.515 95.675 120.885 ;
        RECT 116.330 120.515 117.870 120.885 ;
        RECT 138.525 120.515 140.065 120.885 ;
        RECT 60.845 117.795 62.385 118.165 ;
        RECT 83.040 117.795 84.580 118.165 ;
        RECT 105.235 117.795 106.775 118.165 ;
        RECT 127.430 117.795 128.970 118.165 ;
        RECT 71.940 115.075 73.480 115.445 ;
        RECT 94.135 115.075 95.675 115.445 ;
        RECT 116.330 115.075 117.870 115.445 ;
        RECT 138.525 115.075 140.065 115.445 ;
        RECT 60.845 112.355 62.385 112.725 ;
        RECT 83.040 112.355 84.580 112.725 ;
        RECT 105.235 112.355 106.775 112.725 ;
        RECT 127.430 112.355 128.970 112.725 ;
        RECT 71.940 109.635 73.480 110.005 ;
        RECT 94.135 109.635 95.675 110.005 ;
        RECT 116.330 109.635 117.870 110.005 ;
        RECT 138.525 109.635 140.065 110.005 ;
        RECT 63.960 108.470 64.220 108.790 ;
        RECT 60.845 106.915 62.385 107.285 ;
        RECT 57.060 105.410 57.320 105.730 ;
        RECT 60.280 105.410 60.540 105.730 ;
        RECT 62.580 105.410 62.840 105.730 ;
        RECT 57.120 104.030 57.260 105.410 ;
        RECT 58.900 105.070 59.160 105.390 ;
        RECT 58.960 104.905 59.100 105.070 ;
        RECT 58.890 104.535 59.170 104.905 ;
        RECT 57.060 103.710 57.320 104.030 ;
        RECT 60.340 103.350 60.480 105.410 ;
        RECT 48.780 103.030 49.040 103.350 ;
        RECT 60.280 103.030 60.540 103.350 ;
        RECT 48.840 101.505 48.980 103.030 ;
        RECT 62.640 103.010 62.780 105.410 ;
        RECT 63.500 103.370 63.760 103.690 ;
        RECT 62.580 102.690 62.840 103.010 ;
        RECT 48.770 101.135 49.050 101.505 ;
        RECT 60.845 101.475 62.385 101.845 ;
        RECT 58.900 99.970 59.160 100.290 ;
        RECT 58.440 99.290 58.700 99.610 ;
        RECT 58.500 94.850 58.640 99.290 ;
        RECT 58.960 98.105 59.100 99.970 ;
        RECT 62.640 98.590 62.780 102.690 ;
        RECT 62.580 98.270 62.840 98.590 ;
        RECT 58.890 97.735 59.170 98.105 ;
        RECT 60.280 97.590 60.540 97.910 ;
        RECT 58.440 94.530 58.700 94.850 ;
        RECT 57.980 93.850 58.240 94.170 ;
        RECT 58.040 93.150 58.180 93.850 ;
        RECT 58.500 93.150 58.640 94.530 ;
        RECT 60.340 93.150 60.480 97.590 ;
        RECT 60.845 96.035 62.385 96.405 ;
        RECT 57.980 92.830 58.240 93.150 ;
        RECT 58.440 92.830 58.700 93.150 ;
        RECT 60.280 92.830 60.540 93.150 ;
        RECT 58.500 91.870 58.640 92.830 ;
        RECT 62.580 92.150 62.840 92.470 ;
        RECT 58.500 91.730 59.100 91.870 ;
        RECT 58.960 89.750 59.100 91.730 ;
        RECT 60.280 91.130 60.540 91.450 ;
        RECT 58.900 89.430 59.160 89.750 ;
        RECT 60.340 89.410 60.480 91.130 ;
        RECT 60.845 90.595 62.385 90.965 ;
        RECT 62.640 90.430 62.780 92.150 ;
        RECT 63.560 92.130 63.700 103.370 ;
        RECT 64.020 103.010 64.160 108.470 ;
        RECT 83.040 106.915 84.580 107.285 ;
        RECT 105.235 106.915 106.775 107.285 ;
        RECT 127.430 106.915 128.970 107.285 ;
        RECT 71.940 104.195 73.480 104.565 ;
        RECT 94.135 104.195 95.675 104.565 ;
        RECT 116.330 104.195 117.870 104.565 ;
        RECT 138.525 104.195 140.065 104.565 ;
        RECT 63.960 102.690 64.220 103.010 ;
        RECT 64.020 94.850 64.160 102.690 ;
        RECT 83.040 101.475 84.580 101.845 ;
        RECT 105.235 101.475 106.775 101.845 ;
        RECT 127.430 101.475 128.970 101.845 ;
        RECT 71.940 98.755 73.480 99.125 ;
        RECT 94.135 98.755 95.675 99.125 ;
        RECT 116.330 98.755 117.870 99.125 ;
        RECT 138.525 98.755 140.065 99.125 ;
        RECT 83.040 96.035 84.580 96.405 ;
        RECT 105.235 96.035 106.775 96.405 ;
        RECT 127.430 96.035 128.970 96.405 ;
        RECT 63.960 94.530 64.220 94.850 ;
        RECT 66.260 93.850 66.520 94.170 ;
        RECT 66.320 92.470 66.460 93.850 ;
        RECT 71.940 93.315 73.480 93.685 ;
        RECT 94.135 93.315 95.675 93.685 ;
        RECT 116.330 93.315 117.870 93.685 ;
        RECT 138.525 93.315 140.065 93.685 ;
        RECT 66.260 92.150 66.520 92.470 ;
        RECT 63.500 91.810 63.760 92.130 ;
        RECT 83.040 90.595 84.580 90.965 ;
        RECT 105.235 90.595 106.775 90.965 ;
        RECT 127.430 90.595 128.970 90.965 ;
        RECT 62.580 90.110 62.840 90.430 ;
        RECT 60.280 89.090 60.540 89.410 ;
        RECT 71.940 87.875 73.480 88.245 ;
        RECT 94.135 87.875 95.675 88.245 ;
        RECT 116.330 87.875 117.870 88.245 ;
        RECT 138.525 87.875 140.065 88.245 ;
        RECT 60.845 85.155 62.385 85.525 ;
        RECT 83.040 85.155 84.580 85.525 ;
        RECT 105.235 85.155 106.775 85.525 ;
        RECT 127.430 85.155 128.970 85.525 ;
        RECT 71.940 82.435 73.480 82.805 ;
        RECT 94.135 82.435 95.675 82.805 ;
        RECT 116.330 82.435 117.870 82.805 ;
        RECT 138.525 82.435 140.065 82.805 ;
        RECT 60.845 79.715 62.385 80.085 ;
        RECT 83.040 79.715 84.580 80.085 ;
        RECT 105.235 79.715 106.775 80.085 ;
        RECT 127.430 79.715 128.970 80.085 ;
        RECT 71.940 76.995 73.480 77.365 ;
        RECT 94.135 76.995 95.675 77.365 ;
        RECT 116.330 76.995 117.870 77.365 ;
        RECT 138.525 76.995 140.065 77.365 ;
        RECT 60.845 74.275 62.385 74.645 ;
        RECT 83.040 74.275 84.580 74.645 ;
        RECT 105.235 74.275 106.775 74.645 ;
        RECT 127.430 74.275 128.970 74.645 ;
        RECT 71.940 71.555 73.480 71.925 ;
        RECT 94.135 71.555 95.675 71.925 ;
        RECT 116.330 71.555 117.870 71.925 ;
        RECT 138.525 71.555 140.065 71.925 ;
        RECT 60.845 68.835 62.385 69.205 ;
        RECT 83.040 68.835 84.580 69.205 ;
        RECT 105.235 68.835 106.775 69.205 ;
        RECT 127.430 68.835 128.970 69.205 ;
        RECT 71.940 66.115 73.480 66.485 ;
        RECT 94.135 66.115 95.675 66.485 ;
        RECT 116.330 66.115 117.870 66.485 ;
        RECT 138.525 66.115 140.065 66.485 ;
        RECT 60.845 63.395 62.385 63.765 ;
        RECT 83.040 63.395 84.580 63.765 ;
        RECT 105.235 63.395 106.775 63.765 ;
        RECT 127.430 63.395 128.970 63.765 ;
        RECT 71.940 60.675 73.480 61.045 ;
        RECT 94.135 60.675 95.675 61.045 ;
        RECT 116.330 60.675 117.870 61.045 ;
        RECT 138.525 60.675 140.065 61.045 ;
      LAYER via2 ;
        RECT 71.970 136.880 72.250 137.160 ;
        RECT 72.370 136.880 72.650 137.160 ;
        RECT 72.770 136.880 73.050 137.160 ;
        RECT 73.170 136.880 73.450 137.160 ;
        RECT 94.165 136.880 94.445 137.160 ;
        RECT 94.565 136.880 94.845 137.160 ;
        RECT 94.965 136.880 95.245 137.160 ;
        RECT 95.365 136.880 95.645 137.160 ;
        RECT 116.360 136.880 116.640 137.160 ;
        RECT 116.760 136.880 117.040 137.160 ;
        RECT 117.160 136.880 117.440 137.160 ;
        RECT 117.560 136.880 117.840 137.160 ;
        RECT 138.555 136.880 138.835 137.160 ;
        RECT 138.955 136.880 139.235 137.160 ;
        RECT 139.355 136.880 139.635 137.160 ;
        RECT 139.755 136.880 140.035 137.160 ;
        RECT 60.875 134.160 61.155 134.440 ;
        RECT 61.275 134.160 61.555 134.440 ;
        RECT 61.675 134.160 61.955 134.440 ;
        RECT 62.075 134.160 62.355 134.440 ;
        RECT 83.070 134.160 83.350 134.440 ;
        RECT 83.470 134.160 83.750 134.440 ;
        RECT 83.870 134.160 84.150 134.440 ;
        RECT 84.270 134.160 84.550 134.440 ;
        RECT 105.265 134.160 105.545 134.440 ;
        RECT 105.665 134.160 105.945 134.440 ;
        RECT 106.065 134.160 106.345 134.440 ;
        RECT 106.465 134.160 106.745 134.440 ;
        RECT 127.460 134.160 127.740 134.440 ;
        RECT 127.860 134.160 128.140 134.440 ;
        RECT 128.260 134.160 128.540 134.440 ;
        RECT 128.660 134.160 128.940 134.440 ;
        RECT 71.970 131.440 72.250 131.720 ;
        RECT 72.370 131.440 72.650 131.720 ;
        RECT 72.770 131.440 73.050 131.720 ;
        RECT 73.170 131.440 73.450 131.720 ;
        RECT 94.165 131.440 94.445 131.720 ;
        RECT 94.565 131.440 94.845 131.720 ;
        RECT 94.965 131.440 95.245 131.720 ;
        RECT 95.365 131.440 95.645 131.720 ;
        RECT 116.360 131.440 116.640 131.720 ;
        RECT 116.760 131.440 117.040 131.720 ;
        RECT 117.160 131.440 117.440 131.720 ;
        RECT 117.560 131.440 117.840 131.720 ;
        RECT 138.555 131.440 138.835 131.720 ;
        RECT 138.955 131.440 139.235 131.720 ;
        RECT 139.355 131.440 139.635 131.720 ;
        RECT 139.755 131.440 140.035 131.720 ;
        RECT 60.875 128.720 61.155 129.000 ;
        RECT 61.275 128.720 61.555 129.000 ;
        RECT 61.675 128.720 61.955 129.000 ;
        RECT 62.075 128.720 62.355 129.000 ;
        RECT 83.070 128.720 83.350 129.000 ;
        RECT 83.470 128.720 83.750 129.000 ;
        RECT 83.870 128.720 84.150 129.000 ;
        RECT 84.270 128.720 84.550 129.000 ;
        RECT 105.265 128.720 105.545 129.000 ;
        RECT 105.665 128.720 105.945 129.000 ;
        RECT 106.065 128.720 106.345 129.000 ;
        RECT 106.465 128.720 106.745 129.000 ;
        RECT 127.460 128.720 127.740 129.000 ;
        RECT 127.860 128.720 128.140 129.000 ;
        RECT 128.260 128.720 128.540 129.000 ;
        RECT 128.660 128.720 128.940 129.000 ;
        RECT 71.970 126.000 72.250 126.280 ;
        RECT 72.370 126.000 72.650 126.280 ;
        RECT 72.770 126.000 73.050 126.280 ;
        RECT 73.170 126.000 73.450 126.280 ;
        RECT 94.165 126.000 94.445 126.280 ;
        RECT 94.565 126.000 94.845 126.280 ;
        RECT 94.965 126.000 95.245 126.280 ;
        RECT 95.365 126.000 95.645 126.280 ;
        RECT 116.360 126.000 116.640 126.280 ;
        RECT 116.760 126.000 117.040 126.280 ;
        RECT 117.160 126.000 117.440 126.280 ;
        RECT 117.560 126.000 117.840 126.280 ;
        RECT 138.555 126.000 138.835 126.280 ;
        RECT 138.955 126.000 139.235 126.280 ;
        RECT 139.355 126.000 139.635 126.280 ;
        RECT 139.755 126.000 140.035 126.280 ;
        RECT 60.875 123.280 61.155 123.560 ;
        RECT 61.275 123.280 61.555 123.560 ;
        RECT 61.675 123.280 61.955 123.560 ;
        RECT 62.075 123.280 62.355 123.560 ;
        RECT 83.070 123.280 83.350 123.560 ;
        RECT 83.470 123.280 83.750 123.560 ;
        RECT 83.870 123.280 84.150 123.560 ;
        RECT 84.270 123.280 84.550 123.560 ;
        RECT 105.265 123.280 105.545 123.560 ;
        RECT 105.665 123.280 105.945 123.560 ;
        RECT 106.065 123.280 106.345 123.560 ;
        RECT 106.465 123.280 106.745 123.560 ;
        RECT 127.460 123.280 127.740 123.560 ;
        RECT 127.860 123.280 128.140 123.560 ;
        RECT 128.260 123.280 128.540 123.560 ;
        RECT 128.660 123.280 128.940 123.560 ;
        RECT 71.970 120.560 72.250 120.840 ;
        RECT 72.370 120.560 72.650 120.840 ;
        RECT 72.770 120.560 73.050 120.840 ;
        RECT 73.170 120.560 73.450 120.840 ;
        RECT 94.165 120.560 94.445 120.840 ;
        RECT 94.565 120.560 94.845 120.840 ;
        RECT 94.965 120.560 95.245 120.840 ;
        RECT 95.365 120.560 95.645 120.840 ;
        RECT 116.360 120.560 116.640 120.840 ;
        RECT 116.760 120.560 117.040 120.840 ;
        RECT 117.160 120.560 117.440 120.840 ;
        RECT 117.560 120.560 117.840 120.840 ;
        RECT 138.555 120.560 138.835 120.840 ;
        RECT 138.955 120.560 139.235 120.840 ;
        RECT 139.355 120.560 139.635 120.840 ;
        RECT 139.755 120.560 140.035 120.840 ;
        RECT 60.875 117.840 61.155 118.120 ;
        RECT 61.275 117.840 61.555 118.120 ;
        RECT 61.675 117.840 61.955 118.120 ;
        RECT 62.075 117.840 62.355 118.120 ;
        RECT 83.070 117.840 83.350 118.120 ;
        RECT 83.470 117.840 83.750 118.120 ;
        RECT 83.870 117.840 84.150 118.120 ;
        RECT 84.270 117.840 84.550 118.120 ;
        RECT 105.265 117.840 105.545 118.120 ;
        RECT 105.665 117.840 105.945 118.120 ;
        RECT 106.065 117.840 106.345 118.120 ;
        RECT 106.465 117.840 106.745 118.120 ;
        RECT 127.460 117.840 127.740 118.120 ;
        RECT 127.860 117.840 128.140 118.120 ;
        RECT 128.260 117.840 128.540 118.120 ;
        RECT 128.660 117.840 128.940 118.120 ;
        RECT 71.970 115.120 72.250 115.400 ;
        RECT 72.370 115.120 72.650 115.400 ;
        RECT 72.770 115.120 73.050 115.400 ;
        RECT 73.170 115.120 73.450 115.400 ;
        RECT 94.165 115.120 94.445 115.400 ;
        RECT 94.565 115.120 94.845 115.400 ;
        RECT 94.965 115.120 95.245 115.400 ;
        RECT 95.365 115.120 95.645 115.400 ;
        RECT 116.360 115.120 116.640 115.400 ;
        RECT 116.760 115.120 117.040 115.400 ;
        RECT 117.160 115.120 117.440 115.400 ;
        RECT 117.560 115.120 117.840 115.400 ;
        RECT 138.555 115.120 138.835 115.400 ;
        RECT 138.955 115.120 139.235 115.400 ;
        RECT 139.355 115.120 139.635 115.400 ;
        RECT 139.755 115.120 140.035 115.400 ;
        RECT 60.875 112.400 61.155 112.680 ;
        RECT 61.275 112.400 61.555 112.680 ;
        RECT 61.675 112.400 61.955 112.680 ;
        RECT 62.075 112.400 62.355 112.680 ;
        RECT 83.070 112.400 83.350 112.680 ;
        RECT 83.470 112.400 83.750 112.680 ;
        RECT 83.870 112.400 84.150 112.680 ;
        RECT 84.270 112.400 84.550 112.680 ;
        RECT 105.265 112.400 105.545 112.680 ;
        RECT 105.665 112.400 105.945 112.680 ;
        RECT 106.065 112.400 106.345 112.680 ;
        RECT 106.465 112.400 106.745 112.680 ;
        RECT 127.460 112.400 127.740 112.680 ;
        RECT 127.860 112.400 128.140 112.680 ;
        RECT 128.260 112.400 128.540 112.680 ;
        RECT 128.660 112.400 128.940 112.680 ;
        RECT 71.970 109.680 72.250 109.960 ;
        RECT 72.370 109.680 72.650 109.960 ;
        RECT 72.770 109.680 73.050 109.960 ;
        RECT 73.170 109.680 73.450 109.960 ;
        RECT 94.165 109.680 94.445 109.960 ;
        RECT 94.565 109.680 94.845 109.960 ;
        RECT 94.965 109.680 95.245 109.960 ;
        RECT 95.365 109.680 95.645 109.960 ;
        RECT 116.360 109.680 116.640 109.960 ;
        RECT 116.760 109.680 117.040 109.960 ;
        RECT 117.160 109.680 117.440 109.960 ;
        RECT 117.560 109.680 117.840 109.960 ;
        RECT 138.555 109.680 138.835 109.960 ;
        RECT 138.955 109.680 139.235 109.960 ;
        RECT 139.355 109.680 139.635 109.960 ;
        RECT 139.755 109.680 140.035 109.960 ;
        RECT 60.875 106.960 61.155 107.240 ;
        RECT 61.275 106.960 61.555 107.240 ;
        RECT 61.675 106.960 61.955 107.240 ;
        RECT 62.075 106.960 62.355 107.240 ;
        RECT 58.890 104.580 59.170 104.860 ;
        RECT 60.875 101.520 61.155 101.800 ;
        RECT 61.275 101.520 61.555 101.800 ;
        RECT 61.675 101.520 61.955 101.800 ;
        RECT 62.075 101.520 62.355 101.800 ;
        RECT 48.770 101.180 49.050 101.460 ;
        RECT 58.890 97.780 59.170 98.060 ;
        RECT 60.875 96.080 61.155 96.360 ;
        RECT 61.275 96.080 61.555 96.360 ;
        RECT 61.675 96.080 61.955 96.360 ;
        RECT 62.075 96.080 62.355 96.360 ;
        RECT 60.875 90.640 61.155 90.920 ;
        RECT 61.275 90.640 61.555 90.920 ;
        RECT 61.675 90.640 61.955 90.920 ;
        RECT 62.075 90.640 62.355 90.920 ;
        RECT 83.070 106.960 83.350 107.240 ;
        RECT 83.470 106.960 83.750 107.240 ;
        RECT 83.870 106.960 84.150 107.240 ;
        RECT 84.270 106.960 84.550 107.240 ;
        RECT 105.265 106.960 105.545 107.240 ;
        RECT 105.665 106.960 105.945 107.240 ;
        RECT 106.065 106.960 106.345 107.240 ;
        RECT 106.465 106.960 106.745 107.240 ;
        RECT 127.460 106.960 127.740 107.240 ;
        RECT 127.860 106.960 128.140 107.240 ;
        RECT 128.260 106.960 128.540 107.240 ;
        RECT 128.660 106.960 128.940 107.240 ;
        RECT 71.970 104.240 72.250 104.520 ;
        RECT 72.370 104.240 72.650 104.520 ;
        RECT 72.770 104.240 73.050 104.520 ;
        RECT 73.170 104.240 73.450 104.520 ;
        RECT 94.165 104.240 94.445 104.520 ;
        RECT 94.565 104.240 94.845 104.520 ;
        RECT 94.965 104.240 95.245 104.520 ;
        RECT 95.365 104.240 95.645 104.520 ;
        RECT 116.360 104.240 116.640 104.520 ;
        RECT 116.760 104.240 117.040 104.520 ;
        RECT 117.160 104.240 117.440 104.520 ;
        RECT 117.560 104.240 117.840 104.520 ;
        RECT 138.555 104.240 138.835 104.520 ;
        RECT 138.955 104.240 139.235 104.520 ;
        RECT 139.355 104.240 139.635 104.520 ;
        RECT 139.755 104.240 140.035 104.520 ;
        RECT 83.070 101.520 83.350 101.800 ;
        RECT 83.470 101.520 83.750 101.800 ;
        RECT 83.870 101.520 84.150 101.800 ;
        RECT 84.270 101.520 84.550 101.800 ;
        RECT 105.265 101.520 105.545 101.800 ;
        RECT 105.665 101.520 105.945 101.800 ;
        RECT 106.065 101.520 106.345 101.800 ;
        RECT 106.465 101.520 106.745 101.800 ;
        RECT 127.460 101.520 127.740 101.800 ;
        RECT 127.860 101.520 128.140 101.800 ;
        RECT 128.260 101.520 128.540 101.800 ;
        RECT 128.660 101.520 128.940 101.800 ;
        RECT 71.970 98.800 72.250 99.080 ;
        RECT 72.370 98.800 72.650 99.080 ;
        RECT 72.770 98.800 73.050 99.080 ;
        RECT 73.170 98.800 73.450 99.080 ;
        RECT 94.165 98.800 94.445 99.080 ;
        RECT 94.565 98.800 94.845 99.080 ;
        RECT 94.965 98.800 95.245 99.080 ;
        RECT 95.365 98.800 95.645 99.080 ;
        RECT 116.360 98.800 116.640 99.080 ;
        RECT 116.760 98.800 117.040 99.080 ;
        RECT 117.160 98.800 117.440 99.080 ;
        RECT 117.560 98.800 117.840 99.080 ;
        RECT 138.555 98.800 138.835 99.080 ;
        RECT 138.955 98.800 139.235 99.080 ;
        RECT 139.355 98.800 139.635 99.080 ;
        RECT 139.755 98.800 140.035 99.080 ;
        RECT 83.070 96.080 83.350 96.360 ;
        RECT 83.470 96.080 83.750 96.360 ;
        RECT 83.870 96.080 84.150 96.360 ;
        RECT 84.270 96.080 84.550 96.360 ;
        RECT 105.265 96.080 105.545 96.360 ;
        RECT 105.665 96.080 105.945 96.360 ;
        RECT 106.065 96.080 106.345 96.360 ;
        RECT 106.465 96.080 106.745 96.360 ;
        RECT 127.460 96.080 127.740 96.360 ;
        RECT 127.860 96.080 128.140 96.360 ;
        RECT 128.260 96.080 128.540 96.360 ;
        RECT 128.660 96.080 128.940 96.360 ;
        RECT 71.970 93.360 72.250 93.640 ;
        RECT 72.370 93.360 72.650 93.640 ;
        RECT 72.770 93.360 73.050 93.640 ;
        RECT 73.170 93.360 73.450 93.640 ;
        RECT 94.165 93.360 94.445 93.640 ;
        RECT 94.565 93.360 94.845 93.640 ;
        RECT 94.965 93.360 95.245 93.640 ;
        RECT 95.365 93.360 95.645 93.640 ;
        RECT 116.360 93.360 116.640 93.640 ;
        RECT 116.760 93.360 117.040 93.640 ;
        RECT 117.160 93.360 117.440 93.640 ;
        RECT 117.560 93.360 117.840 93.640 ;
        RECT 138.555 93.360 138.835 93.640 ;
        RECT 138.955 93.360 139.235 93.640 ;
        RECT 139.355 93.360 139.635 93.640 ;
        RECT 139.755 93.360 140.035 93.640 ;
        RECT 83.070 90.640 83.350 90.920 ;
        RECT 83.470 90.640 83.750 90.920 ;
        RECT 83.870 90.640 84.150 90.920 ;
        RECT 84.270 90.640 84.550 90.920 ;
        RECT 105.265 90.640 105.545 90.920 ;
        RECT 105.665 90.640 105.945 90.920 ;
        RECT 106.065 90.640 106.345 90.920 ;
        RECT 106.465 90.640 106.745 90.920 ;
        RECT 127.460 90.640 127.740 90.920 ;
        RECT 127.860 90.640 128.140 90.920 ;
        RECT 128.260 90.640 128.540 90.920 ;
        RECT 128.660 90.640 128.940 90.920 ;
        RECT 71.970 87.920 72.250 88.200 ;
        RECT 72.370 87.920 72.650 88.200 ;
        RECT 72.770 87.920 73.050 88.200 ;
        RECT 73.170 87.920 73.450 88.200 ;
        RECT 94.165 87.920 94.445 88.200 ;
        RECT 94.565 87.920 94.845 88.200 ;
        RECT 94.965 87.920 95.245 88.200 ;
        RECT 95.365 87.920 95.645 88.200 ;
        RECT 116.360 87.920 116.640 88.200 ;
        RECT 116.760 87.920 117.040 88.200 ;
        RECT 117.160 87.920 117.440 88.200 ;
        RECT 117.560 87.920 117.840 88.200 ;
        RECT 138.555 87.920 138.835 88.200 ;
        RECT 138.955 87.920 139.235 88.200 ;
        RECT 139.355 87.920 139.635 88.200 ;
        RECT 139.755 87.920 140.035 88.200 ;
        RECT 60.875 85.200 61.155 85.480 ;
        RECT 61.275 85.200 61.555 85.480 ;
        RECT 61.675 85.200 61.955 85.480 ;
        RECT 62.075 85.200 62.355 85.480 ;
        RECT 83.070 85.200 83.350 85.480 ;
        RECT 83.470 85.200 83.750 85.480 ;
        RECT 83.870 85.200 84.150 85.480 ;
        RECT 84.270 85.200 84.550 85.480 ;
        RECT 105.265 85.200 105.545 85.480 ;
        RECT 105.665 85.200 105.945 85.480 ;
        RECT 106.065 85.200 106.345 85.480 ;
        RECT 106.465 85.200 106.745 85.480 ;
        RECT 127.460 85.200 127.740 85.480 ;
        RECT 127.860 85.200 128.140 85.480 ;
        RECT 128.260 85.200 128.540 85.480 ;
        RECT 128.660 85.200 128.940 85.480 ;
        RECT 71.970 82.480 72.250 82.760 ;
        RECT 72.370 82.480 72.650 82.760 ;
        RECT 72.770 82.480 73.050 82.760 ;
        RECT 73.170 82.480 73.450 82.760 ;
        RECT 94.165 82.480 94.445 82.760 ;
        RECT 94.565 82.480 94.845 82.760 ;
        RECT 94.965 82.480 95.245 82.760 ;
        RECT 95.365 82.480 95.645 82.760 ;
        RECT 116.360 82.480 116.640 82.760 ;
        RECT 116.760 82.480 117.040 82.760 ;
        RECT 117.160 82.480 117.440 82.760 ;
        RECT 117.560 82.480 117.840 82.760 ;
        RECT 138.555 82.480 138.835 82.760 ;
        RECT 138.955 82.480 139.235 82.760 ;
        RECT 139.355 82.480 139.635 82.760 ;
        RECT 139.755 82.480 140.035 82.760 ;
        RECT 60.875 79.760 61.155 80.040 ;
        RECT 61.275 79.760 61.555 80.040 ;
        RECT 61.675 79.760 61.955 80.040 ;
        RECT 62.075 79.760 62.355 80.040 ;
        RECT 83.070 79.760 83.350 80.040 ;
        RECT 83.470 79.760 83.750 80.040 ;
        RECT 83.870 79.760 84.150 80.040 ;
        RECT 84.270 79.760 84.550 80.040 ;
        RECT 105.265 79.760 105.545 80.040 ;
        RECT 105.665 79.760 105.945 80.040 ;
        RECT 106.065 79.760 106.345 80.040 ;
        RECT 106.465 79.760 106.745 80.040 ;
        RECT 127.460 79.760 127.740 80.040 ;
        RECT 127.860 79.760 128.140 80.040 ;
        RECT 128.260 79.760 128.540 80.040 ;
        RECT 128.660 79.760 128.940 80.040 ;
        RECT 71.970 77.040 72.250 77.320 ;
        RECT 72.370 77.040 72.650 77.320 ;
        RECT 72.770 77.040 73.050 77.320 ;
        RECT 73.170 77.040 73.450 77.320 ;
        RECT 94.165 77.040 94.445 77.320 ;
        RECT 94.565 77.040 94.845 77.320 ;
        RECT 94.965 77.040 95.245 77.320 ;
        RECT 95.365 77.040 95.645 77.320 ;
        RECT 116.360 77.040 116.640 77.320 ;
        RECT 116.760 77.040 117.040 77.320 ;
        RECT 117.160 77.040 117.440 77.320 ;
        RECT 117.560 77.040 117.840 77.320 ;
        RECT 138.555 77.040 138.835 77.320 ;
        RECT 138.955 77.040 139.235 77.320 ;
        RECT 139.355 77.040 139.635 77.320 ;
        RECT 139.755 77.040 140.035 77.320 ;
        RECT 60.875 74.320 61.155 74.600 ;
        RECT 61.275 74.320 61.555 74.600 ;
        RECT 61.675 74.320 61.955 74.600 ;
        RECT 62.075 74.320 62.355 74.600 ;
        RECT 83.070 74.320 83.350 74.600 ;
        RECT 83.470 74.320 83.750 74.600 ;
        RECT 83.870 74.320 84.150 74.600 ;
        RECT 84.270 74.320 84.550 74.600 ;
        RECT 105.265 74.320 105.545 74.600 ;
        RECT 105.665 74.320 105.945 74.600 ;
        RECT 106.065 74.320 106.345 74.600 ;
        RECT 106.465 74.320 106.745 74.600 ;
        RECT 127.460 74.320 127.740 74.600 ;
        RECT 127.860 74.320 128.140 74.600 ;
        RECT 128.260 74.320 128.540 74.600 ;
        RECT 128.660 74.320 128.940 74.600 ;
        RECT 71.970 71.600 72.250 71.880 ;
        RECT 72.370 71.600 72.650 71.880 ;
        RECT 72.770 71.600 73.050 71.880 ;
        RECT 73.170 71.600 73.450 71.880 ;
        RECT 94.165 71.600 94.445 71.880 ;
        RECT 94.565 71.600 94.845 71.880 ;
        RECT 94.965 71.600 95.245 71.880 ;
        RECT 95.365 71.600 95.645 71.880 ;
        RECT 116.360 71.600 116.640 71.880 ;
        RECT 116.760 71.600 117.040 71.880 ;
        RECT 117.160 71.600 117.440 71.880 ;
        RECT 117.560 71.600 117.840 71.880 ;
        RECT 138.555 71.600 138.835 71.880 ;
        RECT 138.955 71.600 139.235 71.880 ;
        RECT 139.355 71.600 139.635 71.880 ;
        RECT 139.755 71.600 140.035 71.880 ;
        RECT 60.875 68.880 61.155 69.160 ;
        RECT 61.275 68.880 61.555 69.160 ;
        RECT 61.675 68.880 61.955 69.160 ;
        RECT 62.075 68.880 62.355 69.160 ;
        RECT 83.070 68.880 83.350 69.160 ;
        RECT 83.470 68.880 83.750 69.160 ;
        RECT 83.870 68.880 84.150 69.160 ;
        RECT 84.270 68.880 84.550 69.160 ;
        RECT 105.265 68.880 105.545 69.160 ;
        RECT 105.665 68.880 105.945 69.160 ;
        RECT 106.065 68.880 106.345 69.160 ;
        RECT 106.465 68.880 106.745 69.160 ;
        RECT 127.460 68.880 127.740 69.160 ;
        RECT 127.860 68.880 128.140 69.160 ;
        RECT 128.260 68.880 128.540 69.160 ;
        RECT 128.660 68.880 128.940 69.160 ;
        RECT 71.970 66.160 72.250 66.440 ;
        RECT 72.370 66.160 72.650 66.440 ;
        RECT 72.770 66.160 73.050 66.440 ;
        RECT 73.170 66.160 73.450 66.440 ;
        RECT 94.165 66.160 94.445 66.440 ;
        RECT 94.565 66.160 94.845 66.440 ;
        RECT 94.965 66.160 95.245 66.440 ;
        RECT 95.365 66.160 95.645 66.440 ;
        RECT 116.360 66.160 116.640 66.440 ;
        RECT 116.760 66.160 117.040 66.440 ;
        RECT 117.160 66.160 117.440 66.440 ;
        RECT 117.560 66.160 117.840 66.440 ;
        RECT 138.555 66.160 138.835 66.440 ;
        RECT 138.955 66.160 139.235 66.440 ;
        RECT 139.355 66.160 139.635 66.440 ;
        RECT 139.755 66.160 140.035 66.440 ;
        RECT 60.875 63.440 61.155 63.720 ;
        RECT 61.275 63.440 61.555 63.720 ;
        RECT 61.675 63.440 61.955 63.720 ;
        RECT 62.075 63.440 62.355 63.720 ;
        RECT 83.070 63.440 83.350 63.720 ;
        RECT 83.470 63.440 83.750 63.720 ;
        RECT 83.870 63.440 84.150 63.720 ;
        RECT 84.270 63.440 84.550 63.720 ;
        RECT 105.265 63.440 105.545 63.720 ;
        RECT 105.665 63.440 105.945 63.720 ;
        RECT 106.065 63.440 106.345 63.720 ;
        RECT 106.465 63.440 106.745 63.720 ;
        RECT 127.460 63.440 127.740 63.720 ;
        RECT 127.860 63.440 128.140 63.720 ;
        RECT 128.260 63.440 128.540 63.720 ;
        RECT 128.660 63.440 128.940 63.720 ;
        RECT 71.970 60.720 72.250 61.000 ;
        RECT 72.370 60.720 72.650 61.000 ;
        RECT 72.770 60.720 73.050 61.000 ;
        RECT 73.170 60.720 73.450 61.000 ;
        RECT 94.165 60.720 94.445 61.000 ;
        RECT 94.565 60.720 94.845 61.000 ;
        RECT 94.965 60.720 95.245 61.000 ;
        RECT 95.365 60.720 95.645 61.000 ;
        RECT 116.360 60.720 116.640 61.000 ;
        RECT 116.760 60.720 117.040 61.000 ;
        RECT 117.160 60.720 117.440 61.000 ;
        RECT 117.560 60.720 117.840 61.000 ;
        RECT 138.555 60.720 138.835 61.000 ;
        RECT 138.955 60.720 139.235 61.000 ;
        RECT 139.355 60.720 139.635 61.000 ;
        RECT 139.755 60.720 140.035 61.000 ;
      LAYER met3 ;
        RECT 71.920 136.855 73.500 137.185 ;
        RECT 94.115 136.855 95.695 137.185 ;
        RECT 116.310 136.855 117.890 137.185 ;
        RECT 138.505 136.855 140.085 137.185 ;
        RECT 60.825 134.135 62.405 134.465 ;
        RECT 83.020 134.135 84.600 134.465 ;
        RECT 105.215 134.135 106.795 134.465 ;
        RECT 127.410 134.135 128.990 134.465 ;
        RECT 71.920 131.415 73.500 131.745 ;
        RECT 94.115 131.415 95.695 131.745 ;
        RECT 116.310 131.415 117.890 131.745 ;
        RECT 138.505 131.415 140.085 131.745 ;
        RECT 60.825 128.695 62.405 129.025 ;
        RECT 83.020 128.695 84.600 129.025 ;
        RECT 105.215 128.695 106.795 129.025 ;
        RECT 127.410 128.695 128.990 129.025 ;
        RECT 71.920 125.975 73.500 126.305 ;
        RECT 94.115 125.975 95.695 126.305 ;
        RECT 116.310 125.975 117.890 126.305 ;
        RECT 138.505 125.975 140.085 126.305 ;
        RECT 60.825 123.255 62.405 123.585 ;
        RECT 83.020 123.255 84.600 123.585 ;
        RECT 105.215 123.255 106.795 123.585 ;
        RECT 127.410 123.255 128.990 123.585 ;
        RECT 71.920 120.535 73.500 120.865 ;
        RECT 94.115 120.535 95.695 120.865 ;
        RECT 116.310 120.535 117.890 120.865 ;
        RECT 138.505 120.535 140.085 120.865 ;
        RECT 60.825 117.815 62.405 118.145 ;
        RECT 83.020 117.815 84.600 118.145 ;
        RECT 105.215 117.815 106.795 118.145 ;
        RECT 127.410 117.815 128.990 118.145 ;
        RECT 71.920 115.095 73.500 115.425 ;
        RECT 94.115 115.095 95.695 115.425 ;
        RECT 116.310 115.095 117.890 115.425 ;
        RECT 138.505 115.095 140.085 115.425 ;
        RECT 60.825 112.375 62.405 112.705 ;
        RECT 83.020 112.375 84.600 112.705 ;
        RECT 105.215 112.375 106.795 112.705 ;
        RECT 127.410 112.375 128.990 112.705 ;
        RECT 71.920 109.655 73.500 109.985 ;
        RECT 94.115 109.655 95.695 109.985 ;
        RECT 116.310 109.655 117.890 109.985 ;
        RECT 138.505 109.655 140.085 109.985 ;
        RECT 60.825 106.935 62.405 107.265 ;
        RECT 83.020 106.935 84.600 107.265 ;
        RECT 105.215 106.935 106.795 107.265 ;
        RECT 127.410 106.935 128.990 107.265 ;
        RECT 37.160 105.120 38.060 105.170 ;
        RECT 37.160 105.020 38.720 105.120 ;
        RECT 35.230 104.870 47.000 105.020 ;
        RECT 58.865 104.870 59.195 104.885 ;
        RECT 35.230 104.570 59.195 104.870 ;
        RECT 35.230 104.420 47.000 104.570 ;
        RECT 58.865 104.555 59.195 104.570 ;
        RECT 37.160 104.270 38.720 104.420 ;
        RECT 37.820 104.220 38.720 104.270 ;
        RECT 71.920 104.215 73.500 104.545 ;
        RECT 94.115 104.215 95.695 104.545 ;
        RECT 116.310 104.215 117.890 104.545 ;
        RECT 138.505 104.215 140.085 104.545 ;
        RECT 33.510 101.620 34.470 101.770 ;
        RECT 33.510 101.470 47.000 101.620 ;
        RECT 60.825 101.495 62.405 101.825 ;
        RECT 83.020 101.495 84.600 101.825 ;
        RECT 105.215 101.495 106.795 101.825 ;
        RECT 127.410 101.495 128.990 101.825 ;
        RECT 48.745 101.470 49.075 101.485 ;
        RECT 33.510 101.170 49.075 101.470 ;
        RECT 33.510 101.020 47.000 101.170 ;
        RECT 48.745 101.155 49.075 101.170 ;
        RECT 33.510 100.870 34.470 101.020 ;
        RECT 71.920 98.775 73.500 99.105 ;
        RECT 94.115 98.775 95.695 99.105 ;
        RECT 116.310 98.775 117.890 99.105 ;
        RECT 138.505 98.775 140.085 99.105 ;
        RECT 39.530 98.220 40.490 98.370 ;
        RECT 39.530 98.070 47.000 98.220 ;
        RECT 58.865 98.070 59.195 98.085 ;
        RECT 39.530 97.770 59.195 98.070 ;
        RECT 39.530 97.620 47.000 97.770 ;
        RECT 58.865 97.755 59.195 97.770 ;
        RECT 39.530 97.470 40.490 97.620 ;
        RECT 60.825 96.055 62.405 96.385 ;
        RECT 83.020 96.055 84.600 96.385 ;
        RECT 105.215 96.055 106.795 96.385 ;
        RECT 127.410 96.055 128.990 96.385 ;
        RECT 71.920 93.335 73.500 93.665 ;
        RECT 94.115 93.335 95.695 93.665 ;
        RECT 116.310 93.335 117.890 93.665 ;
        RECT 138.505 93.335 140.085 93.665 ;
        RECT 60.825 90.615 62.405 90.945 ;
        RECT 83.020 90.615 84.600 90.945 ;
        RECT 105.215 90.615 106.795 90.945 ;
        RECT 127.410 90.615 128.990 90.945 ;
        RECT 71.920 87.895 73.500 88.225 ;
        RECT 94.115 87.895 95.695 88.225 ;
        RECT 116.310 87.895 117.890 88.225 ;
        RECT 138.505 87.895 140.085 88.225 ;
        RECT 60.825 85.175 62.405 85.505 ;
        RECT 83.020 85.175 84.600 85.505 ;
        RECT 105.215 85.175 106.795 85.505 ;
        RECT 127.410 85.175 128.990 85.505 ;
        RECT 71.920 82.455 73.500 82.785 ;
        RECT 94.115 82.455 95.695 82.785 ;
        RECT 116.310 82.455 117.890 82.785 ;
        RECT 138.505 82.455 140.085 82.785 ;
        RECT 60.825 79.735 62.405 80.065 ;
        RECT 83.020 79.735 84.600 80.065 ;
        RECT 105.215 79.735 106.795 80.065 ;
        RECT 127.410 79.735 128.990 80.065 ;
        RECT 71.920 77.015 73.500 77.345 ;
        RECT 94.115 77.015 95.695 77.345 ;
        RECT 116.310 77.015 117.890 77.345 ;
        RECT 138.505 77.015 140.085 77.345 ;
        RECT 60.825 74.295 62.405 74.625 ;
        RECT 83.020 74.295 84.600 74.625 ;
        RECT 105.215 74.295 106.795 74.625 ;
        RECT 127.410 74.295 128.990 74.625 ;
        RECT 71.920 71.575 73.500 71.905 ;
        RECT 94.115 71.575 95.695 71.905 ;
        RECT 116.310 71.575 117.890 71.905 ;
        RECT 138.505 71.575 140.085 71.905 ;
        RECT 60.825 68.855 62.405 69.185 ;
        RECT 83.020 68.855 84.600 69.185 ;
        RECT 105.215 68.855 106.795 69.185 ;
        RECT 127.410 68.855 128.990 69.185 ;
        RECT 71.920 66.135 73.500 66.465 ;
        RECT 94.115 66.135 95.695 66.465 ;
        RECT 116.310 66.135 117.890 66.465 ;
        RECT 138.505 66.135 140.085 66.465 ;
        RECT 60.825 63.415 62.405 63.745 ;
        RECT 83.020 63.415 84.600 63.745 ;
        RECT 105.215 63.415 106.795 63.745 ;
        RECT 127.410 63.415 128.990 63.745 ;
        RECT 71.920 60.695 73.500 61.025 ;
        RECT 94.115 60.695 95.695 61.025 ;
        RECT 116.310 60.695 117.890 61.025 ;
        RECT 138.505 60.695 140.085 61.025 ;
      LAYER via3 ;
        RECT 71.950 136.860 72.270 137.180 ;
        RECT 72.350 136.860 72.670 137.180 ;
        RECT 72.750 136.860 73.070 137.180 ;
        RECT 73.150 136.860 73.470 137.180 ;
        RECT 94.145 136.860 94.465 137.180 ;
        RECT 94.545 136.860 94.865 137.180 ;
        RECT 94.945 136.860 95.265 137.180 ;
        RECT 95.345 136.860 95.665 137.180 ;
        RECT 116.340 136.860 116.660 137.180 ;
        RECT 116.740 136.860 117.060 137.180 ;
        RECT 117.140 136.860 117.460 137.180 ;
        RECT 117.540 136.860 117.860 137.180 ;
        RECT 138.535 136.860 138.855 137.180 ;
        RECT 138.935 136.860 139.255 137.180 ;
        RECT 139.335 136.860 139.655 137.180 ;
        RECT 139.735 136.860 140.055 137.180 ;
        RECT 60.855 134.140 61.175 134.460 ;
        RECT 61.255 134.140 61.575 134.460 ;
        RECT 61.655 134.140 61.975 134.460 ;
        RECT 62.055 134.140 62.375 134.460 ;
        RECT 83.050 134.140 83.370 134.460 ;
        RECT 83.450 134.140 83.770 134.460 ;
        RECT 83.850 134.140 84.170 134.460 ;
        RECT 84.250 134.140 84.570 134.460 ;
        RECT 105.245 134.140 105.565 134.460 ;
        RECT 105.645 134.140 105.965 134.460 ;
        RECT 106.045 134.140 106.365 134.460 ;
        RECT 106.445 134.140 106.765 134.460 ;
        RECT 127.440 134.140 127.760 134.460 ;
        RECT 127.840 134.140 128.160 134.460 ;
        RECT 128.240 134.140 128.560 134.460 ;
        RECT 128.640 134.140 128.960 134.460 ;
        RECT 71.950 131.420 72.270 131.740 ;
        RECT 72.350 131.420 72.670 131.740 ;
        RECT 72.750 131.420 73.070 131.740 ;
        RECT 73.150 131.420 73.470 131.740 ;
        RECT 94.145 131.420 94.465 131.740 ;
        RECT 94.545 131.420 94.865 131.740 ;
        RECT 94.945 131.420 95.265 131.740 ;
        RECT 95.345 131.420 95.665 131.740 ;
        RECT 116.340 131.420 116.660 131.740 ;
        RECT 116.740 131.420 117.060 131.740 ;
        RECT 117.140 131.420 117.460 131.740 ;
        RECT 117.540 131.420 117.860 131.740 ;
        RECT 138.535 131.420 138.855 131.740 ;
        RECT 138.935 131.420 139.255 131.740 ;
        RECT 139.335 131.420 139.655 131.740 ;
        RECT 139.735 131.420 140.055 131.740 ;
        RECT 60.855 128.700 61.175 129.020 ;
        RECT 61.255 128.700 61.575 129.020 ;
        RECT 61.655 128.700 61.975 129.020 ;
        RECT 62.055 128.700 62.375 129.020 ;
        RECT 83.050 128.700 83.370 129.020 ;
        RECT 83.450 128.700 83.770 129.020 ;
        RECT 83.850 128.700 84.170 129.020 ;
        RECT 84.250 128.700 84.570 129.020 ;
        RECT 105.245 128.700 105.565 129.020 ;
        RECT 105.645 128.700 105.965 129.020 ;
        RECT 106.045 128.700 106.365 129.020 ;
        RECT 106.445 128.700 106.765 129.020 ;
        RECT 127.440 128.700 127.760 129.020 ;
        RECT 127.840 128.700 128.160 129.020 ;
        RECT 128.240 128.700 128.560 129.020 ;
        RECT 128.640 128.700 128.960 129.020 ;
        RECT 71.950 125.980 72.270 126.300 ;
        RECT 72.350 125.980 72.670 126.300 ;
        RECT 72.750 125.980 73.070 126.300 ;
        RECT 73.150 125.980 73.470 126.300 ;
        RECT 94.145 125.980 94.465 126.300 ;
        RECT 94.545 125.980 94.865 126.300 ;
        RECT 94.945 125.980 95.265 126.300 ;
        RECT 95.345 125.980 95.665 126.300 ;
        RECT 116.340 125.980 116.660 126.300 ;
        RECT 116.740 125.980 117.060 126.300 ;
        RECT 117.140 125.980 117.460 126.300 ;
        RECT 117.540 125.980 117.860 126.300 ;
        RECT 138.535 125.980 138.855 126.300 ;
        RECT 138.935 125.980 139.255 126.300 ;
        RECT 139.335 125.980 139.655 126.300 ;
        RECT 139.735 125.980 140.055 126.300 ;
        RECT 60.855 123.260 61.175 123.580 ;
        RECT 61.255 123.260 61.575 123.580 ;
        RECT 61.655 123.260 61.975 123.580 ;
        RECT 62.055 123.260 62.375 123.580 ;
        RECT 83.050 123.260 83.370 123.580 ;
        RECT 83.450 123.260 83.770 123.580 ;
        RECT 83.850 123.260 84.170 123.580 ;
        RECT 84.250 123.260 84.570 123.580 ;
        RECT 105.245 123.260 105.565 123.580 ;
        RECT 105.645 123.260 105.965 123.580 ;
        RECT 106.045 123.260 106.365 123.580 ;
        RECT 106.445 123.260 106.765 123.580 ;
        RECT 127.440 123.260 127.760 123.580 ;
        RECT 127.840 123.260 128.160 123.580 ;
        RECT 128.240 123.260 128.560 123.580 ;
        RECT 128.640 123.260 128.960 123.580 ;
        RECT 71.950 120.540 72.270 120.860 ;
        RECT 72.350 120.540 72.670 120.860 ;
        RECT 72.750 120.540 73.070 120.860 ;
        RECT 73.150 120.540 73.470 120.860 ;
        RECT 94.145 120.540 94.465 120.860 ;
        RECT 94.545 120.540 94.865 120.860 ;
        RECT 94.945 120.540 95.265 120.860 ;
        RECT 95.345 120.540 95.665 120.860 ;
        RECT 116.340 120.540 116.660 120.860 ;
        RECT 116.740 120.540 117.060 120.860 ;
        RECT 117.140 120.540 117.460 120.860 ;
        RECT 117.540 120.540 117.860 120.860 ;
        RECT 138.535 120.540 138.855 120.860 ;
        RECT 138.935 120.540 139.255 120.860 ;
        RECT 139.335 120.540 139.655 120.860 ;
        RECT 139.735 120.540 140.055 120.860 ;
        RECT 60.855 117.820 61.175 118.140 ;
        RECT 61.255 117.820 61.575 118.140 ;
        RECT 61.655 117.820 61.975 118.140 ;
        RECT 62.055 117.820 62.375 118.140 ;
        RECT 83.050 117.820 83.370 118.140 ;
        RECT 83.450 117.820 83.770 118.140 ;
        RECT 83.850 117.820 84.170 118.140 ;
        RECT 84.250 117.820 84.570 118.140 ;
        RECT 105.245 117.820 105.565 118.140 ;
        RECT 105.645 117.820 105.965 118.140 ;
        RECT 106.045 117.820 106.365 118.140 ;
        RECT 106.445 117.820 106.765 118.140 ;
        RECT 127.440 117.820 127.760 118.140 ;
        RECT 127.840 117.820 128.160 118.140 ;
        RECT 128.240 117.820 128.560 118.140 ;
        RECT 128.640 117.820 128.960 118.140 ;
        RECT 71.950 115.100 72.270 115.420 ;
        RECT 72.350 115.100 72.670 115.420 ;
        RECT 72.750 115.100 73.070 115.420 ;
        RECT 73.150 115.100 73.470 115.420 ;
        RECT 94.145 115.100 94.465 115.420 ;
        RECT 94.545 115.100 94.865 115.420 ;
        RECT 94.945 115.100 95.265 115.420 ;
        RECT 95.345 115.100 95.665 115.420 ;
        RECT 116.340 115.100 116.660 115.420 ;
        RECT 116.740 115.100 117.060 115.420 ;
        RECT 117.140 115.100 117.460 115.420 ;
        RECT 117.540 115.100 117.860 115.420 ;
        RECT 138.535 115.100 138.855 115.420 ;
        RECT 138.935 115.100 139.255 115.420 ;
        RECT 139.335 115.100 139.655 115.420 ;
        RECT 139.735 115.100 140.055 115.420 ;
        RECT 60.855 112.380 61.175 112.700 ;
        RECT 61.255 112.380 61.575 112.700 ;
        RECT 61.655 112.380 61.975 112.700 ;
        RECT 62.055 112.380 62.375 112.700 ;
        RECT 83.050 112.380 83.370 112.700 ;
        RECT 83.450 112.380 83.770 112.700 ;
        RECT 83.850 112.380 84.170 112.700 ;
        RECT 84.250 112.380 84.570 112.700 ;
        RECT 105.245 112.380 105.565 112.700 ;
        RECT 105.645 112.380 105.965 112.700 ;
        RECT 106.045 112.380 106.365 112.700 ;
        RECT 106.445 112.380 106.765 112.700 ;
        RECT 127.440 112.380 127.760 112.700 ;
        RECT 127.840 112.380 128.160 112.700 ;
        RECT 128.240 112.380 128.560 112.700 ;
        RECT 128.640 112.380 128.960 112.700 ;
        RECT 71.950 109.660 72.270 109.980 ;
        RECT 72.350 109.660 72.670 109.980 ;
        RECT 72.750 109.660 73.070 109.980 ;
        RECT 73.150 109.660 73.470 109.980 ;
        RECT 94.145 109.660 94.465 109.980 ;
        RECT 94.545 109.660 94.865 109.980 ;
        RECT 94.945 109.660 95.265 109.980 ;
        RECT 95.345 109.660 95.665 109.980 ;
        RECT 116.340 109.660 116.660 109.980 ;
        RECT 116.740 109.660 117.060 109.980 ;
        RECT 117.140 109.660 117.460 109.980 ;
        RECT 117.540 109.660 117.860 109.980 ;
        RECT 138.535 109.660 138.855 109.980 ;
        RECT 138.935 109.660 139.255 109.980 ;
        RECT 139.335 109.660 139.655 109.980 ;
        RECT 139.735 109.660 140.055 109.980 ;
        RECT 60.855 106.940 61.175 107.260 ;
        RECT 61.255 106.940 61.575 107.260 ;
        RECT 61.655 106.940 61.975 107.260 ;
        RECT 62.055 106.940 62.375 107.260 ;
        RECT 83.050 106.940 83.370 107.260 ;
        RECT 83.450 106.940 83.770 107.260 ;
        RECT 83.850 106.940 84.170 107.260 ;
        RECT 84.250 106.940 84.570 107.260 ;
        RECT 105.245 106.940 105.565 107.260 ;
        RECT 105.645 106.940 105.965 107.260 ;
        RECT 106.045 106.940 106.365 107.260 ;
        RECT 106.445 106.940 106.765 107.260 ;
        RECT 127.440 106.940 127.760 107.260 ;
        RECT 127.840 106.940 128.160 107.260 ;
        RECT 128.240 106.940 128.560 107.260 ;
        RECT 128.640 106.940 128.960 107.260 ;
        RECT 37.250 104.360 37.970 105.080 ;
        RECT 71.950 104.220 72.270 104.540 ;
        RECT 72.350 104.220 72.670 104.540 ;
        RECT 72.750 104.220 73.070 104.540 ;
        RECT 73.150 104.220 73.470 104.540 ;
        RECT 94.145 104.220 94.465 104.540 ;
        RECT 94.545 104.220 94.865 104.540 ;
        RECT 94.945 104.220 95.265 104.540 ;
        RECT 95.345 104.220 95.665 104.540 ;
        RECT 116.340 104.220 116.660 104.540 ;
        RECT 116.740 104.220 117.060 104.540 ;
        RECT 117.140 104.220 117.460 104.540 ;
        RECT 117.540 104.220 117.860 104.540 ;
        RECT 138.535 104.220 138.855 104.540 ;
        RECT 138.935 104.220 139.255 104.540 ;
        RECT 139.335 104.220 139.655 104.540 ;
        RECT 139.735 104.220 140.055 104.540 ;
        RECT 33.630 100.960 34.350 101.680 ;
        RECT 60.855 101.500 61.175 101.820 ;
        RECT 61.255 101.500 61.575 101.820 ;
        RECT 61.655 101.500 61.975 101.820 ;
        RECT 62.055 101.500 62.375 101.820 ;
        RECT 83.050 101.500 83.370 101.820 ;
        RECT 83.450 101.500 83.770 101.820 ;
        RECT 83.850 101.500 84.170 101.820 ;
        RECT 84.250 101.500 84.570 101.820 ;
        RECT 105.245 101.500 105.565 101.820 ;
        RECT 105.645 101.500 105.965 101.820 ;
        RECT 106.045 101.500 106.365 101.820 ;
        RECT 106.445 101.500 106.765 101.820 ;
        RECT 127.440 101.500 127.760 101.820 ;
        RECT 127.840 101.500 128.160 101.820 ;
        RECT 128.240 101.500 128.560 101.820 ;
        RECT 128.640 101.500 128.960 101.820 ;
        RECT 71.950 98.780 72.270 99.100 ;
        RECT 72.350 98.780 72.670 99.100 ;
        RECT 72.750 98.780 73.070 99.100 ;
        RECT 73.150 98.780 73.470 99.100 ;
        RECT 94.145 98.780 94.465 99.100 ;
        RECT 94.545 98.780 94.865 99.100 ;
        RECT 94.945 98.780 95.265 99.100 ;
        RECT 95.345 98.780 95.665 99.100 ;
        RECT 116.340 98.780 116.660 99.100 ;
        RECT 116.740 98.780 117.060 99.100 ;
        RECT 117.140 98.780 117.460 99.100 ;
        RECT 117.540 98.780 117.860 99.100 ;
        RECT 138.535 98.780 138.855 99.100 ;
        RECT 138.935 98.780 139.255 99.100 ;
        RECT 139.335 98.780 139.655 99.100 ;
        RECT 139.735 98.780 140.055 99.100 ;
        RECT 39.650 97.560 40.370 98.280 ;
        RECT 60.855 96.060 61.175 96.380 ;
        RECT 61.255 96.060 61.575 96.380 ;
        RECT 61.655 96.060 61.975 96.380 ;
        RECT 62.055 96.060 62.375 96.380 ;
        RECT 83.050 96.060 83.370 96.380 ;
        RECT 83.450 96.060 83.770 96.380 ;
        RECT 83.850 96.060 84.170 96.380 ;
        RECT 84.250 96.060 84.570 96.380 ;
        RECT 105.245 96.060 105.565 96.380 ;
        RECT 105.645 96.060 105.965 96.380 ;
        RECT 106.045 96.060 106.365 96.380 ;
        RECT 106.445 96.060 106.765 96.380 ;
        RECT 127.440 96.060 127.760 96.380 ;
        RECT 127.840 96.060 128.160 96.380 ;
        RECT 128.240 96.060 128.560 96.380 ;
        RECT 128.640 96.060 128.960 96.380 ;
        RECT 71.950 93.340 72.270 93.660 ;
        RECT 72.350 93.340 72.670 93.660 ;
        RECT 72.750 93.340 73.070 93.660 ;
        RECT 73.150 93.340 73.470 93.660 ;
        RECT 94.145 93.340 94.465 93.660 ;
        RECT 94.545 93.340 94.865 93.660 ;
        RECT 94.945 93.340 95.265 93.660 ;
        RECT 95.345 93.340 95.665 93.660 ;
        RECT 116.340 93.340 116.660 93.660 ;
        RECT 116.740 93.340 117.060 93.660 ;
        RECT 117.140 93.340 117.460 93.660 ;
        RECT 117.540 93.340 117.860 93.660 ;
        RECT 138.535 93.340 138.855 93.660 ;
        RECT 138.935 93.340 139.255 93.660 ;
        RECT 139.335 93.340 139.655 93.660 ;
        RECT 139.735 93.340 140.055 93.660 ;
        RECT 60.855 90.620 61.175 90.940 ;
        RECT 61.255 90.620 61.575 90.940 ;
        RECT 61.655 90.620 61.975 90.940 ;
        RECT 62.055 90.620 62.375 90.940 ;
        RECT 83.050 90.620 83.370 90.940 ;
        RECT 83.450 90.620 83.770 90.940 ;
        RECT 83.850 90.620 84.170 90.940 ;
        RECT 84.250 90.620 84.570 90.940 ;
        RECT 105.245 90.620 105.565 90.940 ;
        RECT 105.645 90.620 105.965 90.940 ;
        RECT 106.045 90.620 106.365 90.940 ;
        RECT 106.445 90.620 106.765 90.940 ;
        RECT 127.440 90.620 127.760 90.940 ;
        RECT 127.840 90.620 128.160 90.940 ;
        RECT 128.240 90.620 128.560 90.940 ;
        RECT 128.640 90.620 128.960 90.940 ;
        RECT 71.950 87.900 72.270 88.220 ;
        RECT 72.350 87.900 72.670 88.220 ;
        RECT 72.750 87.900 73.070 88.220 ;
        RECT 73.150 87.900 73.470 88.220 ;
        RECT 94.145 87.900 94.465 88.220 ;
        RECT 94.545 87.900 94.865 88.220 ;
        RECT 94.945 87.900 95.265 88.220 ;
        RECT 95.345 87.900 95.665 88.220 ;
        RECT 116.340 87.900 116.660 88.220 ;
        RECT 116.740 87.900 117.060 88.220 ;
        RECT 117.140 87.900 117.460 88.220 ;
        RECT 117.540 87.900 117.860 88.220 ;
        RECT 138.535 87.900 138.855 88.220 ;
        RECT 138.935 87.900 139.255 88.220 ;
        RECT 139.335 87.900 139.655 88.220 ;
        RECT 139.735 87.900 140.055 88.220 ;
        RECT 60.855 85.180 61.175 85.500 ;
        RECT 61.255 85.180 61.575 85.500 ;
        RECT 61.655 85.180 61.975 85.500 ;
        RECT 62.055 85.180 62.375 85.500 ;
        RECT 83.050 85.180 83.370 85.500 ;
        RECT 83.450 85.180 83.770 85.500 ;
        RECT 83.850 85.180 84.170 85.500 ;
        RECT 84.250 85.180 84.570 85.500 ;
        RECT 105.245 85.180 105.565 85.500 ;
        RECT 105.645 85.180 105.965 85.500 ;
        RECT 106.045 85.180 106.365 85.500 ;
        RECT 106.445 85.180 106.765 85.500 ;
        RECT 127.440 85.180 127.760 85.500 ;
        RECT 127.840 85.180 128.160 85.500 ;
        RECT 128.240 85.180 128.560 85.500 ;
        RECT 128.640 85.180 128.960 85.500 ;
        RECT 71.950 82.460 72.270 82.780 ;
        RECT 72.350 82.460 72.670 82.780 ;
        RECT 72.750 82.460 73.070 82.780 ;
        RECT 73.150 82.460 73.470 82.780 ;
        RECT 94.145 82.460 94.465 82.780 ;
        RECT 94.545 82.460 94.865 82.780 ;
        RECT 94.945 82.460 95.265 82.780 ;
        RECT 95.345 82.460 95.665 82.780 ;
        RECT 116.340 82.460 116.660 82.780 ;
        RECT 116.740 82.460 117.060 82.780 ;
        RECT 117.140 82.460 117.460 82.780 ;
        RECT 117.540 82.460 117.860 82.780 ;
        RECT 138.535 82.460 138.855 82.780 ;
        RECT 138.935 82.460 139.255 82.780 ;
        RECT 139.335 82.460 139.655 82.780 ;
        RECT 139.735 82.460 140.055 82.780 ;
        RECT 60.855 79.740 61.175 80.060 ;
        RECT 61.255 79.740 61.575 80.060 ;
        RECT 61.655 79.740 61.975 80.060 ;
        RECT 62.055 79.740 62.375 80.060 ;
        RECT 83.050 79.740 83.370 80.060 ;
        RECT 83.450 79.740 83.770 80.060 ;
        RECT 83.850 79.740 84.170 80.060 ;
        RECT 84.250 79.740 84.570 80.060 ;
        RECT 105.245 79.740 105.565 80.060 ;
        RECT 105.645 79.740 105.965 80.060 ;
        RECT 106.045 79.740 106.365 80.060 ;
        RECT 106.445 79.740 106.765 80.060 ;
        RECT 127.440 79.740 127.760 80.060 ;
        RECT 127.840 79.740 128.160 80.060 ;
        RECT 128.240 79.740 128.560 80.060 ;
        RECT 128.640 79.740 128.960 80.060 ;
        RECT 71.950 77.020 72.270 77.340 ;
        RECT 72.350 77.020 72.670 77.340 ;
        RECT 72.750 77.020 73.070 77.340 ;
        RECT 73.150 77.020 73.470 77.340 ;
        RECT 94.145 77.020 94.465 77.340 ;
        RECT 94.545 77.020 94.865 77.340 ;
        RECT 94.945 77.020 95.265 77.340 ;
        RECT 95.345 77.020 95.665 77.340 ;
        RECT 116.340 77.020 116.660 77.340 ;
        RECT 116.740 77.020 117.060 77.340 ;
        RECT 117.140 77.020 117.460 77.340 ;
        RECT 117.540 77.020 117.860 77.340 ;
        RECT 138.535 77.020 138.855 77.340 ;
        RECT 138.935 77.020 139.255 77.340 ;
        RECT 139.335 77.020 139.655 77.340 ;
        RECT 139.735 77.020 140.055 77.340 ;
        RECT 60.855 74.300 61.175 74.620 ;
        RECT 61.255 74.300 61.575 74.620 ;
        RECT 61.655 74.300 61.975 74.620 ;
        RECT 62.055 74.300 62.375 74.620 ;
        RECT 83.050 74.300 83.370 74.620 ;
        RECT 83.450 74.300 83.770 74.620 ;
        RECT 83.850 74.300 84.170 74.620 ;
        RECT 84.250 74.300 84.570 74.620 ;
        RECT 105.245 74.300 105.565 74.620 ;
        RECT 105.645 74.300 105.965 74.620 ;
        RECT 106.045 74.300 106.365 74.620 ;
        RECT 106.445 74.300 106.765 74.620 ;
        RECT 127.440 74.300 127.760 74.620 ;
        RECT 127.840 74.300 128.160 74.620 ;
        RECT 128.240 74.300 128.560 74.620 ;
        RECT 128.640 74.300 128.960 74.620 ;
        RECT 71.950 71.580 72.270 71.900 ;
        RECT 72.350 71.580 72.670 71.900 ;
        RECT 72.750 71.580 73.070 71.900 ;
        RECT 73.150 71.580 73.470 71.900 ;
        RECT 94.145 71.580 94.465 71.900 ;
        RECT 94.545 71.580 94.865 71.900 ;
        RECT 94.945 71.580 95.265 71.900 ;
        RECT 95.345 71.580 95.665 71.900 ;
        RECT 116.340 71.580 116.660 71.900 ;
        RECT 116.740 71.580 117.060 71.900 ;
        RECT 117.140 71.580 117.460 71.900 ;
        RECT 117.540 71.580 117.860 71.900 ;
        RECT 138.535 71.580 138.855 71.900 ;
        RECT 138.935 71.580 139.255 71.900 ;
        RECT 139.335 71.580 139.655 71.900 ;
        RECT 139.735 71.580 140.055 71.900 ;
        RECT 60.855 68.860 61.175 69.180 ;
        RECT 61.255 68.860 61.575 69.180 ;
        RECT 61.655 68.860 61.975 69.180 ;
        RECT 62.055 68.860 62.375 69.180 ;
        RECT 83.050 68.860 83.370 69.180 ;
        RECT 83.450 68.860 83.770 69.180 ;
        RECT 83.850 68.860 84.170 69.180 ;
        RECT 84.250 68.860 84.570 69.180 ;
        RECT 105.245 68.860 105.565 69.180 ;
        RECT 105.645 68.860 105.965 69.180 ;
        RECT 106.045 68.860 106.365 69.180 ;
        RECT 106.445 68.860 106.765 69.180 ;
        RECT 127.440 68.860 127.760 69.180 ;
        RECT 127.840 68.860 128.160 69.180 ;
        RECT 128.240 68.860 128.560 69.180 ;
        RECT 128.640 68.860 128.960 69.180 ;
        RECT 71.950 66.140 72.270 66.460 ;
        RECT 72.350 66.140 72.670 66.460 ;
        RECT 72.750 66.140 73.070 66.460 ;
        RECT 73.150 66.140 73.470 66.460 ;
        RECT 94.145 66.140 94.465 66.460 ;
        RECT 94.545 66.140 94.865 66.460 ;
        RECT 94.945 66.140 95.265 66.460 ;
        RECT 95.345 66.140 95.665 66.460 ;
        RECT 116.340 66.140 116.660 66.460 ;
        RECT 116.740 66.140 117.060 66.460 ;
        RECT 117.140 66.140 117.460 66.460 ;
        RECT 117.540 66.140 117.860 66.460 ;
        RECT 138.535 66.140 138.855 66.460 ;
        RECT 138.935 66.140 139.255 66.460 ;
        RECT 139.335 66.140 139.655 66.460 ;
        RECT 139.735 66.140 140.055 66.460 ;
        RECT 60.855 63.420 61.175 63.740 ;
        RECT 61.255 63.420 61.575 63.740 ;
        RECT 61.655 63.420 61.975 63.740 ;
        RECT 62.055 63.420 62.375 63.740 ;
        RECT 83.050 63.420 83.370 63.740 ;
        RECT 83.450 63.420 83.770 63.740 ;
        RECT 83.850 63.420 84.170 63.740 ;
        RECT 84.250 63.420 84.570 63.740 ;
        RECT 105.245 63.420 105.565 63.740 ;
        RECT 105.645 63.420 105.965 63.740 ;
        RECT 106.045 63.420 106.365 63.740 ;
        RECT 106.445 63.420 106.765 63.740 ;
        RECT 127.440 63.420 127.760 63.740 ;
        RECT 127.840 63.420 128.160 63.740 ;
        RECT 128.240 63.420 128.560 63.740 ;
        RECT 128.640 63.420 128.960 63.740 ;
        RECT 71.950 60.700 72.270 61.020 ;
        RECT 72.350 60.700 72.670 61.020 ;
        RECT 72.750 60.700 73.070 61.020 ;
        RECT 73.150 60.700 73.470 61.020 ;
        RECT 94.145 60.700 94.465 61.020 ;
        RECT 94.545 60.700 94.865 61.020 ;
        RECT 94.945 60.700 95.265 61.020 ;
        RECT 95.345 60.700 95.665 61.020 ;
        RECT 116.340 60.700 116.660 61.020 ;
        RECT 116.740 60.700 117.060 61.020 ;
        RECT 117.140 60.700 117.460 61.020 ;
        RECT 117.540 60.700 117.860 61.020 ;
        RECT 138.535 60.700 138.855 61.020 ;
        RECT 138.935 60.700 139.255 61.020 ;
        RECT 139.335 60.700 139.655 61.020 ;
        RECT 139.735 60.700 140.055 61.020 ;
      LAYER met4 ;
        RECT 6.000 4.980 8.000 220.740 ;
        RECT 9.000 220.450 11.000 220.740 ;
        RECT 35.670 220.450 35.970 225.740 ;
        RECT 38.430 220.450 38.730 225.740 ;
        RECT 41.190 220.450 41.490 225.740 ;
        RECT 43.950 220.450 44.250 225.740 ;
        RECT 46.710 220.450 47.010 225.740 ;
        RECT 49.470 220.450 49.770 225.740 ;
        RECT 52.230 220.450 52.530 225.740 ;
        RECT 54.990 220.450 55.290 225.740 ;
        RECT 57.750 220.450 58.050 225.740 ;
        RECT 60.510 220.450 60.810 225.740 ;
        RECT 63.270 220.450 63.570 225.740 ;
        RECT 66.030 220.450 66.330 225.740 ;
        RECT 68.790 220.450 69.090 225.740 ;
        RECT 71.550 220.450 71.850 225.740 ;
        RECT 74.310 220.450 74.610 225.740 ;
        RECT 77.070 220.450 77.370 225.740 ;
        RECT 79.830 224.740 80.130 225.740 ;
        RECT 82.590 224.740 82.890 225.740 ;
        RECT 85.350 224.740 85.650 225.740 ;
        RECT 88.110 224.740 88.410 225.740 ;
        RECT 90.870 224.740 91.170 225.740 ;
        RECT 93.630 224.740 93.930 225.740 ;
        RECT 96.390 224.740 96.690 225.740 ;
        RECT 99.150 224.740 99.450 225.740 ;
        RECT 101.910 224.740 102.210 225.740 ;
        RECT 104.670 224.740 104.970 225.740 ;
        RECT 107.430 224.740 107.730 225.740 ;
        RECT 110.190 224.740 110.490 225.740 ;
        RECT 112.950 224.740 113.250 225.740 ;
        RECT 115.710 224.740 116.010 225.740 ;
        RECT 118.470 224.740 118.770 225.740 ;
        RECT 121.230 224.740 121.530 225.740 ;
        RECT 123.990 224.740 124.290 225.740 ;
        RECT 126.750 224.740 127.050 225.740 ;
        RECT 129.510 224.740 129.810 225.740 ;
        RECT 132.270 224.740 132.570 225.740 ;
        RECT 135.030 224.740 135.330 225.740 ;
        RECT 137.790 224.740 138.090 225.740 ;
        RECT 140.550 224.740 140.850 225.740 ;
        RECT 143.310 224.740 143.610 225.740 ;
        RECT 146.070 224.740 146.370 225.740 ;
        RECT 148.830 224.740 149.130 225.740 ;
        RECT 151.590 224.740 151.890 225.740 ;
        RECT 9.000 218.450 86.820 220.450 ;
        RECT 9.000 4.980 11.000 218.450 ;
        RECT 32.800 161.450 157.710 162.350 ;
        RECT 32.800 105.120 33.700 161.450 ;
        RECT 37.155 105.120 38.065 105.175 ;
        RECT 32.800 104.220 38.720 105.120 ;
        RECT 33.535 101.770 34.445 101.775 ;
        RECT 28.700 100.870 38.660 101.770 ;
        RECT 28.700 42.860 29.600 100.870 ;
        RECT 33.535 100.865 34.445 100.870 ;
        RECT 39.555 98.350 40.465 98.375 ;
        RECT 37.690 97.450 42.110 98.350 ;
        RECT 37.690 51.240 38.590 97.450 ;
        RECT 60.815 60.620 62.415 137.260 ;
        RECT 71.910 60.620 73.510 137.260 ;
        RECT 83.010 60.620 84.610 137.260 ;
        RECT 94.105 60.620 95.705 137.260 ;
        RECT 105.205 60.620 106.805 137.260 ;
        RECT 116.300 60.620 117.900 137.260 ;
        RECT 127.400 60.620 129.000 137.260 ;
        RECT 138.495 60.620 140.095 137.260 ;
        RECT 37.690 50.340 138.390 51.240 ;
        RECT 28.700 41.960 119.070 42.860 ;
        RECT 21.570 -0.020 22.470 0.980 ;
        RECT 40.890 -0.020 41.790 0.980 ;
        RECT 60.210 -0.020 61.110 0.980 ;
        RECT 79.530 -0.020 80.430 0.980 ;
        RECT 98.850 -0.020 99.750 0.980 ;
        RECT 118.170 -0.020 119.070 41.960 ;
        RECT 137.490 -0.020 138.390 50.340 ;
        RECT 156.810 -0.020 157.710 161.450 ;
  END
END tt_um_brandonramos_opamp_ladder
END LIBRARY

