VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test_1
  CLASS BLOCK ;
  FOREIGN tt_um_test_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.601000 ;
    PORT
      LAYER met3 ;
        RECT 159.000 108.840 161.000 109.440 ;
    END
  END Out
  PIN VGND
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.910 10.640 61.510 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.780 10.640 100.380 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.650 10.640 139.250 215.120 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 40.475 10.640 42.075 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.345 10.640 80.945 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.215 10.640 119.815 215.120 ;
    END
  END VPWR
  PIN Vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 159.000 115.640 161.000 116.240 ;
    END
  END Vin
  PIN Vip
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 159.000 112.240 161.000 112.840 ;
    END
  END Vip
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 155.670 215.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 155.480 214.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 155.480 215.120 ;
      LAYER met2 ;
        RECT 21.070 10.695 154.010 215.065 ;
      LAYER met3 ;
        RECT 21.050 116.640 159.000 215.045 ;
        RECT 21.050 115.240 158.600 116.640 ;
        RECT 21.050 113.240 159.000 115.240 ;
        RECT 21.050 111.840 158.600 113.240 ;
        RECT 21.050 109.840 159.000 111.840 ;
        RECT 21.050 108.440 158.600 109.840 ;
        RECT 21.050 10.715 159.000 108.440 ;
  END
END tt_um_test_1
END LIBRARY

