VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_brandonramos_opamp_ladder
  CLASS BLOCK ;
  FOREIGN tt_um_brandonramos_opamp_ladder ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  OBS
      LAYER pwell ;
        RECT 50.665 136.925 50.835 137.095 ;
        RECT 52.045 136.925 52.215 137.095 ;
        RECT 57.565 136.925 57.735 137.095 ;
        RECT 63.080 136.955 63.200 137.065 ;
        RECT 64.005 136.925 64.175 137.095 ;
        RECT 69.525 136.925 69.695 137.095 ;
        RECT 75.045 136.925 75.215 137.095 ;
        RECT 76.885 136.925 77.055 137.095 ;
        RECT 82.405 136.925 82.575 137.095 ;
        RECT 87.925 136.925 88.095 137.095 ;
        RECT 89.765 136.925 89.935 137.095 ;
        RECT 95.285 136.925 95.455 137.095 ;
        RECT 100.805 136.925 100.975 137.095 ;
        RECT 102.645 136.925 102.815 137.095 ;
        RECT 108.165 136.925 108.335 137.095 ;
        RECT 113.685 136.925 113.855 137.095 ;
        RECT 115.525 136.925 115.695 137.095 ;
        RECT 121.045 136.925 121.215 137.095 ;
        RECT 126.565 136.925 126.735 137.095 ;
        RECT 128.405 136.925 128.575 137.095 ;
        RECT 133.925 136.925 134.095 137.095 ;
        RECT 137.600 136.955 137.720 137.065 ;
        RECT 138.985 136.925 139.155 137.095 ;
        RECT 63.545 136.165 63.715 136.690 ;
        RECT 76.425 136.165 76.595 136.690 ;
        RECT 89.305 136.165 89.475 136.690 ;
        RECT 102.185 136.165 102.355 136.690 ;
        RECT 115.065 136.165 115.235 136.690 ;
        RECT 127.945 136.165 128.115 136.690 ;
      LAYER nwell ;
        RECT 50.330 132.875 139.490 135.705 ;
      LAYER pwell ;
        RECT 63.545 131.890 63.715 132.415 ;
        RECT 89.305 131.890 89.475 132.415 ;
        RECT 115.065 131.890 115.235 132.415 ;
        RECT 50.665 131.485 50.835 131.655 ;
        RECT 52.045 131.485 52.215 131.655 ;
        RECT 57.565 131.485 57.735 131.655 ;
        RECT 63.085 131.625 63.255 131.655 ;
        RECT 63.080 131.515 63.255 131.625 ;
        RECT 63.085 131.485 63.255 131.515 ;
        RECT 64.005 131.485 64.175 131.655 ;
        RECT 68.605 131.485 68.775 131.655 ;
        RECT 69.525 131.485 69.695 131.655 ;
        RECT 74.125 131.485 74.295 131.655 ;
        RECT 75.045 131.485 75.215 131.655 ;
        RECT 75.960 131.515 76.080 131.625 ;
        RECT 76.885 131.485 77.055 131.655 ;
        RECT 80.565 131.485 80.735 131.655 ;
        RECT 82.405 131.485 82.575 131.655 ;
        RECT 86.085 131.485 86.255 131.655 ;
        RECT 87.925 131.485 88.095 131.655 ;
        RECT 88.840 131.515 88.960 131.625 ;
        RECT 89.765 131.485 89.935 131.655 ;
        RECT 93.445 131.485 93.615 131.655 ;
        RECT 95.285 131.485 95.455 131.655 ;
        RECT 98.965 131.485 99.135 131.655 ;
        RECT 100.805 131.485 100.975 131.655 ;
        RECT 101.720 131.515 101.840 131.625 ;
        RECT 102.645 131.485 102.815 131.655 ;
        RECT 106.325 131.485 106.495 131.655 ;
        RECT 108.165 131.485 108.335 131.655 ;
        RECT 111.845 131.485 112.015 131.655 ;
        RECT 113.685 131.485 113.855 131.655 ;
        RECT 114.600 131.515 114.720 131.625 ;
        RECT 115.525 131.485 115.695 131.655 ;
        RECT 119.205 131.485 119.375 131.655 ;
        RECT 121.045 131.485 121.215 131.655 ;
        RECT 124.725 131.485 124.895 131.655 ;
        RECT 126.565 131.485 126.735 131.655 ;
        RECT 127.480 131.515 127.600 131.625 ;
        RECT 128.405 131.485 128.575 131.655 ;
        RECT 132.085 131.485 132.255 131.655 ;
        RECT 133.925 131.485 134.095 131.655 ;
        RECT 137.600 131.515 137.720 131.625 ;
        RECT 138.985 131.485 139.155 131.655 ;
        RECT 76.425 130.725 76.595 131.250 ;
        RECT 102.185 130.725 102.355 131.250 ;
        RECT 127.945 130.725 128.115 131.250 ;
      LAYER nwell ;
        RECT 50.330 127.435 139.490 130.265 ;
      LAYER pwell ;
        RECT 63.545 126.450 63.715 126.975 ;
        RECT 89.305 126.450 89.475 126.975 ;
        RECT 115.065 126.450 115.235 126.975 ;
        RECT 50.665 126.045 50.835 126.215 ;
        RECT 52.045 126.045 52.215 126.215 ;
        RECT 57.565 126.045 57.735 126.215 ;
        RECT 63.085 126.185 63.255 126.215 ;
        RECT 63.080 126.075 63.255 126.185 ;
        RECT 63.085 126.045 63.255 126.075 ;
        RECT 64.005 126.045 64.175 126.215 ;
        RECT 68.605 126.045 68.775 126.215 ;
        RECT 69.525 126.045 69.695 126.215 ;
        RECT 74.125 126.045 74.295 126.215 ;
        RECT 75.045 126.045 75.215 126.215 ;
        RECT 75.960 126.075 76.080 126.185 ;
        RECT 76.885 126.045 77.055 126.215 ;
        RECT 80.565 126.045 80.735 126.215 ;
        RECT 82.405 126.045 82.575 126.215 ;
        RECT 86.085 126.045 86.255 126.215 ;
        RECT 87.925 126.045 88.095 126.215 ;
        RECT 88.840 126.075 88.960 126.185 ;
        RECT 89.765 126.045 89.935 126.215 ;
        RECT 93.445 126.045 93.615 126.215 ;
        RECT 95.285 126.045 95.455 126.215 ;
        RECT 98.965 126.045 99.135 126.215 ;
        RECT 100.805 126.045 100.975 126.215 ;
        RECT 101.720 126.075 101.840 126.185 ;
        RECT 102.645 126.045 102.815 126.215 ;
        RECT 106.325 126.045 106.495 126.215 ;
        RECT 108.165 126.045 108.335 126.215 ;
        RECT 111.845 126.045 112.015 126.215 ;
        RECT 113.685 126.045 113.855 126.215 ;
        RECT 114.600 126.075 114.720 126.185 ;
        RECT 115.525 126.045 115.695 126.215 ;
        RECT 119.205 126.045 119.375 126.215 ;
        RECT 121.045 126.045 121.215 126.215 ;
        RECT 124.725 126.045 124.895 126.215 ;
        RECT 126.565 126.045 126.735 126.215 ;
        RECT 127.480 126.075 127.600 126.185 ;
        RECT 128.405 126.045 128.575 126.215 ;
        RECT 132.085 126.045 132.255 126.215 ;
        RECT 133.925 126.045 134.095 126.215 ;
        RECT 137.600 126.075 137.720 126.185 ;
        RECT 138.985 126.045 139.155 126.215 ;
        RECT 76.425 125.285 76.595 125.810 ;
        RECT 102.185 125.285 102.355 125.810 ;
        RECT 127.945 125.285 128.115 125.810 ;
      LAYER nwell ;
        RECT 50.330 121.995 139.490 124.825 ;
      LAYER pwell ;
        RECT 63.545 121.010 63.715 121.535 ;
        RECT 89.305 121.010 89.475 121.535 ;
        RECT 115.065 121.010 115.235 121.535 ;
        RECT 50.665 120.605 50.835 120.775 ;
        RECT 52.045 120.605 52.215 120.775 ;
        RECT 57.565 120.605 57.735 120.775 ;
        RECT 63.085 120.745 63.255 120.775 ;
        RECT 63.080 120.635 63.255 120.745 ;
        RECT 63.085 120.605 63.255 120.635 ;
        RECT 64.005 120.605 64.175 120.775 ;
        RECT 68.605 120.605 68.775 120.775 ;
        RECT 69.525 120.605 69.695 120.775 ;
        RECT 74.125 120.605 74.295 120.775 ;
        RECT 75.045 120.605 75.215 120.775 ;
        RECT 75.960 120.635 76.080 120.745 ;
        RECT 76.885 120.605 77.055 120.775 ;
        RECT 80.565 120.605 80.735 120.775 ;
        RECT 82.405 120.605 82.575 120.775 ;
        RECT 86.085 120.605 86.255 120.775 ;
        RECT 87.925 120.605 88.095 120.775 ;
        RECT 88.840 120.635 88.960 120.745 ;
        RECT 89.765 120.605 89.935 120.775 ;
        RECT 93.445 120.605 93.615 120.775 ;
        RECT 95.285 120.605 95.455 120.775 ;
        RECT 98.965 120.605 99.135 120.775 ;
        RECT 100.805 120.605 100.975 120.775 ;
        RECT 101.720 120.635 101.840 120.745 ;
        RECT 102.645 120.605 102.815 120.775 ;
        RECT 106.325 120.605 106.495 120.775 ;
        RECT 108.165 120.605 108.335 120.775 ;
        RECT 111.845 120.605 112.015 120.775 ;
        RECT 113.685 120.605 113.855 120.775 ;
        RECT 114.600 120.635 114.720 120.745 ;
        RECT 115.525 120.605 115.695 120.775 ;
        RECT 119.205 120.605 119.375 120.775 ;
        RECT 121.045 120.605 121.215 120.775 ;
        RECT 124.725 120.605 124.895 120.775 ;
        RECT 126.565 120.605 126.735 120.775 ;
        RECT 127.480 120.635 127.600 120.745 ;
        RECT 128.405 120.605 128.575 120.775 ;
        RECT 132.085 120.605 132.255 120.775 ;
        RECT 133.925 120.605 134.095 120.775 ;
        RECT 137.600 120.635 137.720 120.745 ;
        RECT 138.985 120.605 139.155 120.775 ;
        RECT 76.425 119.845 76.595 120.370 ;
        RECT 102.185 119.845 102.355 120.370 ;
        RECT 127.945 119.845 128.115 120.370 ;
      LAYER nwell ;
        RECT 50.330 116.555 139.490 119.385 ;
      LAYER pwell ;
        RECT 63.545 115.570 63.715 116.095 ;
        RECT 89.305 115.570 89.475 116.095 ;
        RECT 115.065 115.570 115.235 116.095 ;
        RECT 50.665 115.165 50.835 115.335 ;
        RECT 52.045 115.165 52.215 115.335 ;
        RECT 57.565 115.165 57.735 115.335 ;
        RECT 63.085 115.305 63.255 115.335 ;
        RECT 63.080 115.195 63.255 115.305 ;
        RECT 63.085 115.165 63.255 115.195 ;
        RECT 64.005 115.165 64.175 115.335 ;
        RECT 68.605 115.165 68.775 115.335 ;
        RECT 69.525 115.165 69.695 115.335 ;
        RECT 74.125 115.165 74.295 115.335 ;
        RECT 75.045 115.165 75.215 115.335 ;
        RECT 75.960 115.195 76.080 115.305 ;
        RECT 76.885 115.165 77.055 115.335 ;
        RECT 80.565 115.165 80.735 115.335 ;
        RECT 82.405 115.165 82.575 115.335 ;
        RECT 86.085 115.165 86.255 115.335 ;
        RECT 87.925 115.165 88.095 115.335 ;
        RECT 88.840 115.195 88.960 115.305 ;
        RECT 89.765 115.165 89.935 115.335 ;
        RECT 93.445 115.165 93.615 115.335 ;
        RECT 95.285 115.165 95.455 115.335 ;
        RECT 98.965 115.165 99.135 115.335 ;
        RECT 100.805 115.165 100.975 115.335 ;
        RECT 101.720 115.195 101.840 115.305 ;
        RECT 102.645 115.165 102.815 115.335 ;
        RECT 106.325 115.165 106.495 115.335 ;
        RECT 108.165 115.165 108.335 115.335 ;
        RECT 111.845 115.165 112.015 115.335 ;
        RECT 113.685 115.165 113.855 115.335 ;
        RECT 114.600 115.195 114.720 115.305 ;
        RECT 115.525 115.165 115.695 115.335 ;
        RECT 119.205 115.165 119.375 115.335 ;
        RECT 121.045 115.165 121.215 115.335 ;
        RECT 124.725 115.165 124.895 115.335 ;
        RECT 126.565 115.165 126.735 115.335 ;
        RECT 127.480 115.195 127.600 115.305 ;
        RECT 128.405 115.165 128.575 115.335 ;
        RECT 132.085 115.165 132.255 115.335 ;
        RECT 133.925 115.165 134.095 115.335 ;
        RECT 137.600 115.195 137.720 115.305 ;
        RECT 138.985 115.165 139.155 115.335 ;
        RECT 76.425 114.405 76.595 114.930 ;
        RECT 102.185 114.405 102.355 114.930 ;
        RECT 127.945 114.405 128.115 114.930 ;
      LAYER nwell ;
        RECT 50.330 111.115 139.490 113.945 ;
      LAYER pwell ;
        RECT 63.545 110.130 63.715 110.655 ;
        RECT 89.305 110.130 89.475 110.655 ;
        RECT 115.065 110.130 115.235 110.655 ;
        RECT 50.665 109.725 50.835 109.895 ;
        RECT 52.045 109.725 52.215 109.895 ;
        RECT 57.565 109.725 57.735 109.895 ;
        RECT 63.085 109.865 63.255 109.895 ;
        RECT 63.080 109.755 63.255 109.865 ;
        RECT 63.085 109.725 63.255 109.755 ;
        RECT 64.005 109.725 64.175 109.895 ;
        RECT 64.920 109.755 65.040 109.865 ;
        RECT 65.385 109.725 65.555 109.895 ;
        RECT 66.765 109.725 66.935 109.895 ;
        RECT 68.605 109.725 68.775 109.895 ;
        RECT 69.525 109.725 69.695 109.895 ;
        RECT 74.125 109.725 74.295 109.895 ;
        RECT 75.045 109.725 75.215 109.895 ;
        RECT 75.960 109.755 76.080 109.865 ;
        RECT 76.885 109.725 77.055 109.895 ;
        RECT 80.565 109.725 80.735 109.895 ;
        RECT 82.405 109.725 82.575 109.895 ;
        RECT 86.085 109.725 86.255 109.895 ;
        RECT 87.925 109.725 88.095 109.895 ;
        RECT 88.840 109.755 88.960 109.865 ;
        RECT 89.765 109.725 89.935 109.895 ;
        RECT 93.445 109.725 93.615 109.895 ;
        RECT 95.285 109.725 95.455 109.895 ;
        RECT 98.965 109.725 99.135 109.895 ;
        RECT 100.805 109.725 100.975 109.895 ;
        RECT 101.720 109.755 101.840 109.865 ;
        RECT 102.645 109.725 102.815 109.895 ;
        RECT 106.325 109.725 106.495 109.895 ;
        RECT 108.165 109.725 108.335 109.895 ;
        RECT 111.845 109.725 112.015 109.895 ;
        RECT 113.685 109.725 113.855 109.895 ;
        RECT 114.600 109.755 114.720 109.865 ;
        RECT 115.525 109.725 115.695 109.895 ;
        RECT 119.205 109.725 119.375 109.895 ;
        RECT 121.045 109.725 121.215 109.895 ;
        RECT 124.725 109.725 124.895 109.895 ;
        RECT 126.565 109.725 126.735 109.895 ;
        RECT 127.480 109.755 127.600 109.865 ;
        RECT 128.405 109.725 128.575 109.895 ;
        RECT 132.085 109.725 132.255 109.895 ;
        RECT 133.925 109.725 134.095 109.895 ;
        RECT 137.600 109.755 137.720 109.865 ;
        RECT 138.985 109.725 139.155 109.895 ;
        RECT 76.425 108.965 76.595 109.490 ;
        RECT 102.185 108.965 102.355 109.490 ;
        RECT 127.945 108.965 128.115 109.490 ;
      LAYER nwell ;
        RECT 50.330 105.675 139.490 108.505 ;
      LAYER pwell ;
        RECT 63.545 104.690 63.715 105.215 ;
        RECT 89.305 104.690 89.475 105.215 ;
        RECT 115.065 104.690 115.235 105.215 ;
        RECT 50.665 104.285 50.835 104.455 ;
        RECT 52.045 104.285 52.225 104.455 ;
        RECT 53.425 104.285 53.595 104.455 ;
        RECT 55.720 104.315 55.840 104.425 ;
        RECT 57.105 104.285 57.275 104.455 ;
        RECT 57.560 104.285 57.730 104.455 ;
        RECT 58.955 104.310 59.115 104.420 ;
        RECT 59.870 104.285 60.040 104.455 ;
        RECT 62.160 104.285 62.340 104.455 ;
        RECT 62.635 104.320 62.795 104.430 ;
        RECT 64.005 104.285 64.175 104.455 ;
        RECT 66.305 104.285 66.475 104.455 ;
        RECT 69.525 104.285 69.695 104.455 ;
        RECT 71.825 104.285 71.995 104.455 ;
        RECT 75.045 104.285 75.215 104.455 ;
        RECT 75.515 104.310 75.675 104.420 ;
        RECT 76.885 104.285 77.055 104.455 ;
        RECT 80.565 104.285 80.735 104.455 ;
        RECT 82.405 104.285 82.575 104.455 ;
        RECT 86.085 104.285 86.255 104.455 ;
        RECT 87.925 104.285 88.095 104.455 ;
        RECT 88.840 104.315 88.960 104.425 ;
        RECT 89.765 104.285 89.935 104.455 ;
        RECT 93.445 104.285 93.615 104.455 ;
        RECT 95.285 104.285 95.455 104.455 ;
        RECT 98.965 104.285 99.135 104.455 ;
        RECT 100.805 104.285 100.975 104.455 ;
        RECT 101.720 104.315 101.840 104.425 ;
        RECT 102.645 104.285 102.815 104.455 ;
        RECT 106.325 104.285 106.495 104.455 ;
        RECT 108.165 104.285 108.335 104.455 ;
        RECT 111.845 104.285 112.015 104.455 ;
        RECT 113.685 104.285 113.855 104.455 ;
        RECT 114.600 104.315 114.720 104.425 ;
        RECT 115.525 104.285 115.695 104.455 ;
        RECT 119.205 104.285 119.375 104.455 ;
        RECT 121.045 104.285 121.215 104.455 ;
        RECT 124.725 104.285 124.895 104.455 ;
        RECT 126.565 104.285 126.735 104.455 ;
        RECT 127.480 104.315 127.600 104.425 ;
        RECT 128.405 104.285 128.575 104.455 ;
        RECT 132.085 104.285 132.255 104.455 ;
        RECT 133.925 104.285 134.095 104.455 ;
        RECT 137.600 104.315 137.720 104.425 ;
        RECT 138.985 104.285 139.155 104.455 ;
        RECT 76.425 103.525 76.595 104.050 ;
        RECT 102.185 103.525 102.355 104.050 ;
        RECT 127.945 103.525 128.115 104.050 ;
      LAYER nwell ;
        RECT 50.330 100.235 139.490 103.065 ;
      LAYER pwell ;
        RECT 63.545 99.250 63.715 99.775 ;
        RECT 89.305 99.250 89.475 99.775 ;
        RECT 115.065 99.250 115.235 99.775 ;
        RECT 50.665 98.845 50.835 99.015 ;
        RECT 52.045 98.845 52.225 99.015 ;
        RECT 53.425 98.845 53.595 99.015 ;
        RECT 57.565 98.845 57.735 99.015 ;
        RECT 58.945 98.845 59.115 99.015 ;
        RECT 60.320 98.875 60.440 98.985 ;
        RECT 60.785 98.845 60.955 99.015 ;
        RECT 62.165 98.845 62.335 99.015 ;
        RECT 62.635 98.880 62.795 98.990 ;
        RECT 64.005 98.845 64.175 99.015 ;
        RECT 67.685 98.845 67.855 99.015 ;
        RECT 69.525 98.845 69.695 99.015 ;
        RECT 73.205 98.845 73.375 99.015 ;
        RECT 75.045 98.845 75.215 99.015 ;
        RECT 75.960 98.875 76.080 98.985 ;
        RECT 76.885 98.845 77.055 99.015 ;
        RECT 80.565 98.845 80.735 99.015 ;
        RECT 82.405 98.845 82.575 99.015 ;
        RECT 86.085 98.845 86.255 99.015 ;
        RECT 87.925 98.845 88.095 99.015 ;
        RECT 88.840 98.875 88.960 98.985 ;
        RECT 89.765 98.845 89.935 99.015 ;
        RECT 93.445 98.845 93.615 99.015 ;
        RECT 95.285 98.845 95.455 99.015 ;
        RECT 98.965 98.845 99.135 99.015 ;
        RECT 100.805 98.845 100.975 99.015 ;
        RECT 101.720 98.875 101.840 98.985 ;
        RECT 102.645 98.845 102.815 99.015 ;
        RECT 106.325 98.845 106.495 99.015 ;
        RECT 108.165 98.845 108.335 99.015 ;
        RECT 111.845 98.845 112.015 99.015 ;
        RECT 113.685 98.845 113.855 99.015 ;
        RECT 114.600 98.875 114.720 98.985 ;
        RECT 115.525 98.845 115.695 99.015 ;
        RECT 119.205 98.845 119.375 99.015 ;
        RECT 121.045 98.845 121.215 99.015 ;
        RECT 124.725 98.845 124.895 99.015 ;
        RECT 126.565 98.845 126.735 99.015 ;
        RECT 127.480 98.875 127.600 98.985 ;
        RECT 128.405 98.845 128.575 99.015 ;
        RECT 132.085 98.845 132.255 99.015 ;
        RECT 133.925 98.845 134.095 99.015 ;
        RECT 137.600 98.875 137.720 98.985 ;
        RECT 138.985 98.845 139.155 99.015 ;
        RECT 76.425 98.085 76.595 98.610 ;
        RECT 102.185 98.085 102.355 98.610 ;
        RECT 127.945 98.085 128.115 98.610 ;
      LAYER nwell ;
        RECT 50.330 94.795 139.490 97.625 ;
      LAYER pwell ;
        RECT 63.545 93.810 63.715 94.335 ;
        RECT 89.305 93.810 89.475 94.335 ;
        RECT 115.065 93.810 115.235 94.335 ;
        RECT 50.665 93.405 50.835 93.575 ;
        RECT 52.045 93.405 52.215 93.575 ;
        RECT 55.735 93.430 55.895 93.540 ;
        RECT 57.565 93.405 57.735 93.575 ;
        RECT 60.050 93.405 60.220 93.575 ;
        RECT 61.060 93.405 61.230 93.575 ;
        RECT 61.240 93.435 61.360 93.545 ;
        RECT 62.630 93.405 62.800 93.575 ;
        RECT 63.080 93.435 63.200 93.545 ;
        RECT 64.005 93.405 64.175 93.575 ;
        RECT 64.925 93.405 65.095 93.575 ;
        RECT 66.305 93.405 66.475 93.575 ;
        RECT 67.685 93.405 67.855 93.575 ;
        RECT 69.525 93.405 69.695 93.575 ;
        RECT 73.205 93.405 73.375 93.575 ;
        RECT 75.045 93.405 75.215 93.575 ;
        RECT 75.960 93.435 76.080 93.545 ;
        RECT 76.885 93.405 77.055 93.575 ;
        RECT 80.565 93.405 80.735 93.575 ;
        RECT 82.405 93.405 82.575 93.575 ;
        RECT 86.085 93.405 86.255 93.575 ;
        RECT 87.925 93.405 88.095 93.575 ;
        RECT 88.840 93.435 88.960 93.545 ;
        RECT 89.765 93.405 89.935 93.575 ;
        RECT 93.445 93.405 93.615 93.575 ;
        RECT 95.285 93.405 95.455 93.575 ;
        RECT 98.965 93.405 99.135 93.575 ;
        RECT 100.805 93.405 100.975 93.575 ;
        RECT 101.720 93.435 101.840 93.545 ;
        RECT 102.645 93.405 102.815 93.575 ;
        RECT 106.325 93.405 106.495 93.575 ;
        RECT 108.165 93.405 108.335 93.575 ;
        RECT 111.845 93.405 112.015 93.575 ;
        RECT 113.685 93.405 113.855 93.575 ;
        RECT 114.600 93.435 114.720 93.545 ;
        RECT 115.525 93.405 115.695 93.575 ;
        RECT 119.205 93.405 119.375 93.575 ;
        RECT 121.045 93.405 121.215 93.575 ;
        RECT 124.725 93.405 124.895 93.575 ;
        RECT 126.565 93.405 126.735 93.575 ;
        RECT 127.480 93.435 127.600 93.545 ;
        RECT 128.405 93.405 128.575 93.575 ;
        RECT 132.085 93.405 132.255 93.575 ;
        RECT 133.925 93.405 134.095 93.575 ;
        RECT 137.600 93.435 137.720 93.545 ;
        RECT 138.985 93.405 139.155 93.575 ;
        RECT 76.425 92.645 76.595 93.170 ;
        RECT 102.185 92.645 102.355 93.170 ;
        RECT 127.945 92.645 128.115 93.170 ;
      LAYER nwell ;
        RECT 50.330 89.355 139.490 92.185 ;
      LAYER pwell ;
        RECT 63.545 88.370 63.715 88.895 ;
        RECT 89.305 88.370 89.475 88.895 ;
        RECT 115.065 88.370 115.235 88.895 ;
        RECT 50.665 87.965 50.835 88.135 ;
        RECT 52.045 87.965 52.215 88.135 ;
        RECT 57.565 87.965 57.735 88.135 ;
        RECT 60.335 87.965 60.505 88.135 ;
        RECT 61.705 87.965 61.875 88.135 ;
        RECT 63.085 88.105 63.255 88.135 ;
        RECT 63.080 87.995 63.255 88.105 ;
        RECT 63.085 87.965 63.255 87.995 ;
        RECT 64.005 87.965 64.175 88.135 ;
        RECT 68.605 87.965 68.775 88.135 ;
        RECT 69.525 87.965 69.695 88.135 ;
        RECT 74.125 87.965 74.295 88.135 ;
        RECT 75.045 87.965 75.215 88.135 ;
        RECT 75.960 87.995 76.080 88.105 ;
        RECT 76.885 87.965 77.055 88.135 ;
        RECT 80.565 87.965 80.735 88.135 ;
        RECT 82.405 87.965 82.575 88.135 ;
        RECT 86.085 87.965 86.255 88.135 ;
        RECT 87.925 87.965 88.095 88.135 ;
        RECT 88.840 87.995 88.960 88.105 ;
        RECT 89.765 87.965 89.935 88.135 ;
        RECT 93.445 87.965 93.615 88.135 ;
        RECT 95.285 87.965 95.455 88.135 ;
        RECT 98.965 87.965 99.135 88.135 ;
        RECT 100.805 87.965 100.975 88.135 ;
        RECT 101.720 87.995 101.840 88.105 ;
        RECT 102.645 87.965 102.815 88.135 ;
        RECT 106.325 87.965 106.495 88.135 ;
        RECT 108.165 87.965 108.335 88.135 ;
        RECT 111.845 87.965 112.015 88.135 ;
        RECT 113.685 87.965 113.855 88.135 ;
        RECT 114.600 87.995 114.720 88.105 ;
        RECT 115.525 87.965 115.695 88.135 ;
        RECT 119.205 87.965 119.375 88.135 ;
        RECT 121.045 87.965 121.215 88.135 ;
        RECT 124.725 87.965 124.895 88.135 ;
        RECT 126.565 87.965 126.735 88.135 ;
        RECT 127.480 87.995 127.600 88.105 ;
        RECT 128.405 87.965 128.575 88.135 ;
        RECT 132.085 87.965 132.255 88.135 ;
        RECT 133.925 87.965 134.095 88.135 ;
        RECT 137.600 87.995 137.720 88.105 ;
        RECT 138.985 87.965 139.155 88.135 ;
        RECT 76.425 87.205 76.595 87.730 ;
        RECT 102.185 87.205 102.355 87.730 ;
        RECT 127.945 87.205 128.115 87.730 ;
      LAYER nwell ;
        RECT 50.330 83.915 139.490 86.745 ;
      LAYER pwell ;
        RECT 63.545 82.930 63.715 83.455 ;
        RECT 89.305 82.930 89.475 83.455 ;
        RECT 115.065 82.930 115.235 83.455 ;
        RECT 50.665 82.525 50.835 82.695 ;
        RECT 52.045 82.525 52.215 82.695 ;
        RECT 57.565 82.525 57.735 82.695 ;
        RECT 63.085 82.665 63.255 82.695 ;
        RECT 63.080 82.555 63.255 82.665 ;
        RECT 63.085 82.525 63.255 82.555 ;
        RECT 64.005 82.525 64.175 82.695 ;
        RECT 68.605 82.525 68.775 82.695 ;
        RECT 69.525 82.525 69.695 82.695 ;
        RECT 74.125 82.525 74.295 82.695 ;
        RECT 75.045 82.525 75.215 82.695 ;
        RECT 75.960 82.555 76.080 82.665 ;
        RECT 76.885 82.525 77.055 82.695 ;
        RECT 80.565 82.525 80.735 82.695 ;
        RECT 82.405 82.525 82.575 82.695 ;
        RECT 86.085 82.525 86.255 82.695 ;
        RECT 87.925 82.525 88.095 82.695 ;
        RECT 88.840 82.555 88.960 82.665 ;
        RECT 89.765 82.525 89.935 82.695 ;
        RECT 93.445 82.525 93.615 82.695 ;
        RECT 95.285 82.525 95.455 82.695 ;
        RECT 98.965 82.525 99.135 82.695 ;
        RECT 100.805 82.525 100.975 82.695 ;
        RECT 101.720 82.555 101.840 82.665 ;
        RECT 102.645 82.525 102.815 82.695 ;
        RECT 106.325 82.525 106.495 82.695 ;
        RECT 108.165 82.525 108.335 82.695 ;
        RECT 111.845 82.525 112.015 82.695 ;
        RECT 113.685 82.525 113.855 82.695 ;
        RECT 114.600 82.555 114.720 82.665 ;
        RECT 115.525 82.525 115.695 82.695 ;
        RECT 119.205 82.525 119.375 82.695 ;
        RECT 121.045 82.525 121.215 82.695 ;
        RECT 124.725 82.525 124.895 82.695 ;
        RECT 126.565 82.525 126.735 82.695 ;
        RECT 127.480 82.555 127.600 82.665 ;
        RECT 128.405 82.525 128.575 82.695 ;
        RECT 132.085 82.525 132.255 82.695 ;
        RECT 133.925 82.525 134.095 82.695 ;
        RECT 137.600 82.555 137.720 82.665 ;
        RECT 138.985 82.525 139.155 82.695 ;
        RECT 76.425 81.765 76.595 82.290 ;
        RECT 102.185 81.765 102.355 82.290 ;
        RECT 127.945 81.765 128.115 82.290 ;
      LAYER nwell ;
        RECT 50.330 78.475 139.490 81.305 ;
      LAYER pwell ;
        RECT 63.545 77.490 63.715 78.015 ;
        RECT 89.305 77.490 89.475 78.015 ;
        RECT 115.065 77.490 115.235 78.015 ;
        RECT 50.665 77.085 50.835 77.255 ;
        RECT 52.045 77.085 52.215 77.255 ;
        RECT 57.565 77.085 57.735 77.255 ;
        RECT 63.085 77.225 63.255 77.255 ;
        RECT 63.080 77.115 63.255 77.225 ;
        RECT 63.085 77.085 63.255 77.115 ;
        RECT 64.005 77.085 64.175 77.255 ;
        RECT 68.605 77.085 68.775 77.255 ;
        RECT 69.525 77.085 69.695 77.255 ;
        RECT 74.125 77.085 74.295 77.255 ;
        RECT 75.045 77.085 75.215 77.255 ;
        RECT 75.960 77.115 76.080 77.225 ;
        RECT 76.885 77.085 77.055 77.255 ;
        RECT 80.565 77.085 80.735 77.255 ;
        RECT 82.405 77.085 82.575 77.255 ;
        RECT 86.085 77.085 86.255 77.255 ;
        RECT 87.925 77.085 88.095 77.255 ;
        RECT 88.840 77.115 88.960 77.225 ;
        RECT 89.765 77.085 89.935 77.255 ;
        RECT 93.445 77.085 93.615 77.255 ;
        RECT 95.285 77.085 95.455 77.255 ;
        RECT 98.965 77.085 99.135 77.255 ;
        RECT 100.805 77.085 100.975 77.255 ;
        RECT 101.720 77.115 101.840 77.225 ;
        RECT 102.645 77.085 102.815 77.255 ;
        RECT 106.325 77.085 106.495 77.255 ;
        RECT 108.165 77.085 108.335 77.255 ;
        RECT 111.845 77.085 112.015 77.255 ;
        RECT 113.685 77.085 113.855 77.255 ;
        RECT 114.600 77.115 114.720 77.225 ;
        RECT 115.525 77.085 115.695 77.255 ;
        RECT 119.205 77.085 119.375 77.255 ;
        RECT 121.045 77.085 121.215 77.255 ;
        RECT 124.725 77.085 124.895 77.255 ;
        RECT 126.565 77.085 126.735 77.255 ;
        RECT 127.480 77.115 127.600 77.225 ;
        RECT 128.405 77.085 128.575 77.255 ;
        RECT 132.085 77.085 132.255 77.255 ;
        RECT 133.925 77.085 134.095 77.255 ;
        RECT 137.600 77.115 137.720 77.225 ;
        RECT 138.985 77.085 139.155 77.255 ;
        RECT 76.425 76.325 76.595 76.850 ;
        RECT 102.185 76.325 102.355 76.850 ;
        RECT 127.945 76.325 128.115 76.850 ;
      LAYER nwell ;
        RECT 50.330 73.035 139.490 75.865 ;
      LAYER pwell ;
        RECT 63.545 72.050 63.715 72.575 ;
        RECT 89.305 72.050 89.475 72.575 ;
        RECT 115.065 72.050 115.235 72.575 ;
        RECT 50.665 71.645 50.835 71.815 ;
        RECT 52.045 71.645 52.215 71.815 ;
        RECT 57.565 71.645 57.735 71.815 ;
        RECT 63.085 71.785 63.255 71.815 ;
        RECT 63.080 71.675 63.255 71.785 ;
        RECT 63.085 71.645 63.255 71.675 ;
        RECT 64.005 71.645 64.175 71.815 ;
        RECT 68.605 71.645 68.775 71.815 ;
        RECT 69.525 71.645 69.695 71.815 ;
        RECT 74.125 71.645 74.295 71.815 ;
        RECT 75.045 71.645 75.215 71.815 ;
        RECT 75.960 71.675 76.080 71.785 ;
        RECT 76.885 71.645 77.055 71.815 ;
        RECT 80.565 71.645 80.735 71.815 ;
        RECT 82.405 71.645 82.575 71.815 ;
        RECT 86.085 71.645 86.255 71.815 ;
        RECT 87.925 71.645 88.095 71.815 ;
        RECT 88.840 71.675 88.960 71.785 ;
        RECT 89.765 71.645 89.935 71.815 ;
        RECT 93.445 71.645 93.615 71.815 ;
        RECT 95.285 71.645 95.455 71.815 ;
        RECT 98.965 71.645 99.135 71.815 ;
        RECT 100.805 71.645 100.975 71.815 ;
        RECT 101.720 71.675 101.840 71.785 ;
        RECT 102.645 71.645 102.815 71.815 ;
        RECT 106.325 71.645 106.495 71.815 ;
        RECT 108.165 71.645 108.335 71.815 ;
        RECT 111.845 71.645 112.015 71.815 ;
        RECT 113.685 71.645 113.855 71.815 ;
        RECT 114.600 71.675 114.720 71.785 ;
        RECT 115.525 71.645 115.695 71.815 ;
        RECT 119.205 71.645 119.375 71.815 ;
        RECT 121.045 71.645 121.215 71.815 ;
        RECT 124.725 71.645 124.895 71.815 ;
        RECT 126.565 71.645 126.735 71.815 ;
        RECT 127.480 71.675 127.600 71.785 ;
        RECT 128.405 71.645 128.575 71.815 ;
        RECT 132.085 71.645 132.255 71.815 ;
        RECT 133.925 71.645 134.095 71.815 ;
        RECT 137.600 71.675 137.720 71.785 ;
        RECT 138.985 71.645 139.155 71.815 ;
        RECT 76.425 70.885 76.595 71.410 ;
        RECT 102.185 70.885 102.355 71.410 ;
        RECT 127.945 70.885 128.115 71.410 ;
      LAYER nwell ;
        RECT 50.330 67.595 139.490 70.425 ;
      LAYER pwell ;
        RECT 63.545 66.610 63.715 67.135 ;
        RECT 89.305 66.610 89.475 67.135 ;
        RECT 115.065 66.610 115.235 67.135 ;
        RECT 50.665 66.205 50.835 66.375 ;
        RECT 52.045 66.205 52.215 66.375 ;
        RECT 57.565 66.205 57.735 66.375 ;
        RECT 63.085 66.345 63.255 66.375 ;
        RECT 63.080 66.235 63.255 66.345 ;
        RECT 63.085 66.205 63.255 66.235 ;
        RECT 64.005 66.205 64.175 66.375 ;
        RECT 68.605 66.205 68.775 66.375 ;
        RECT 69.525 66.205 69.695 66.375 ;
        RECT 74.125 66.205 74.295 66.375 ;
        RECT 75.045 66.205 75.215 66.375 ;
        RECT 75.960 66.235 76.080 66.345 ;
        RECT 76.885 66.205 77.055 66.375 ;
        RECT 80.565 66.205 80.735 66.375 ;
        RECT 82.405 66.205 82.575 66.375 ;
        RECT 86.085 66.205 86.255 66.375 ;
        RECT 87.925 66.205 88.095 66.375 ;
        RECT 88.840 66.235 88.960 66.345 ;
        RECT 89.765 66.205 89.935 66.375 ;
        RECT 93.445 66.205 93.615 66.375 ;
        RECT 95.285 66.205 95.455 66.375 ;
        RECT 98.965 66.205 99.135 66.375 ;
        RECT 100.805 66.205 100.975 66.375 ;
        RECT 101.720 66.235 101.840 66.345 ;
        RECT 102.645 66.205 102.815 66.375 ;
        RECT 106.325 66.205 106.495 66.375 ;
        RECT 108.165 66.205 108.335 66.375 ;
        RECT 111.845 66.205 112.015 66.375 ;
        RECT 113.685 66.205 113.855 66.375 ;
        RECT 114.600 66.235 114.720 66.345 ;
        RECT 115.525 66.205 115.695 66.375 ;
        RECT 119.205 66.205 119.375 66.375 ;
        RECT 121.045 66.205 121.215 66.375 ;
        RECT 124.725 66.205 124.895 66.375 ;
        RECT 126.565 66.205 126.735 66.375 ;
        RECT 127.480 66.235 127.600 66.345 ;
        RECT 128.405 66.205 128.575 66.375 ;
        RECT 132.085 66.205 132.255 66.375 ;
        RECT 133.925 66.205 134.095 66.375 ;
        RECT 137.600 66.235 137.720 66.345 ;
        RECT 138.985 66.205 139.155 66.375 ;
        RECT 76.425 65.445 76.595 65.970 ;
        RECT 102.185 65.445 102.355 65.970 ;
        RECT 127.945 65.445 128.115 65.970 ;
      LAYER nwell ;
        RECT 50.330 62.155 139.490 64.985 ;
      LAYER pwell ;
        RECT 63.545 61.170 63.715 61.695 ;
        RECT 76.425 61.170 76.595 61.695 ;
        RECT 89.305 61.170 89.475 61.695 ;
        RECT 102.185 61.170 102.355 61.695 ;
        RECT 115.065 61.170 115.235 61.695 ;
        RECT 127.945 61.170 128.115 61.695 ;
        RECT 50.665 60.765 50.835 60.935 ;
        RECT 52.045 60.765 52.215 60.935 ;
        RECT 57.565 60.765 57.735 60.935 ;
        RECT 63.080 60.795 63.200 60.905 ;
        RECT 64.005 60.765 64.175 60.935 ;
        RECT 69.525 60.765 69.695 60.935 ;
        RECT 75.045 60.765 75.215 60.935 ;
        RECT 76.885 60.765 77.055 60.935 ;
        RECT 82.405 60.765 82.575 60.935 ;
        RECT 87.925 60.765 88.095 60.935 ;
        RECT 89.765 60.765 89.935 60.935 ;
        RECT 95.285 60.765 95.455 60.935 ;
        RECT 100.805 60.765 100.975 60.935 ;
        RECT 102.645 60.765 102.815 60.935 ;
        RECT 108.165 60.765 108.335 60.935 ;
        RECT 113.685 60.765 113.855 60.935 ;
        RECT 115.525 60.765 115.695 60.935 ;
        RECT 121.045 60.765 121.215 60.935 ;
        RECT 126.565 60.765 126.735 60.935 ;
        RECT 128.405 60.765 128.575 60.935 ;
        RECT 133.925 60.765 134.095 60.935 ;
        RECT 137.600 60.795 137.720 60.905 ;
        RECT 138.985 60.765 139.155 60.935 ;
      LAYER li1 ;
        RECT 50.520 136.925 139.300 137.095 ;
        RECT 50.605 136.175 51.815 136.925 ;
        RECT 51.985 136.380 57.330 136.925 ;
        RECT 57.505 136.380 62.850 136.925 ;
        RECT 50.605 135.635 51.125 136.175 ;
        RECT 51.295 135.465 51.815 136.005 ;
        RECT 53.570 135.550 53.910 136.380 ;
        RECT 50.605 134.375 51.815 135.465 ;
        RECT 55.390 134.810 55.740 136.060 ;
        RECT 59.090 135.550 59.430 136.380 ;
        RECT 63.485 136.200 63.775 136.925 ;
        RECT 63.945 136.380 69.290 136.925 ;
        RECT 69.465 136.380 74.810 136.925 ;
        RECT 60.910 134.810 61.260 136.060 ;
        RECT 65.530 135.550 65.870 136.380 ;
        RECT 51.985 134.375 57.330 134.810 ;
        RECT 57.505 134.375 62.850 134.810 ;
        RECT 63.485 134.375 63.775 135.540 ;
        RECT 67.350 134.810 67.700 136.060 ;
        RECT 71.050 135.550 71.390 136.380 ;
        RECT 74.985 136.175 76.195 136.925 ;
        RECT 76.365 136.200 76.655 136.925 ;
        RECT 76.825 136.380 82.170 136.925 ;
        RECT 82.345 136.380 87.690 136.925 ;
        RECT 72.870 134.810 73.220 136.060 ;
        RECT 74.985 135.635 75.505 136.175 ;
        RECT 75.675 135.465 76.195 136.005 ;
        RECT 78.410 135.550 78.750 136.380 ;
        RECT 63.945 134.375 69.290 134.810 ;
        RECT 69.465 134.375 74.810 134.810 ;
        RECT 74.985 134.375 76.195 135.465 ;
        RECT 76.365 134.375 76.655 135.540 ;
        RECT 80.230 134.810 80.580 136.060 ;
        RECT 83.930 135.550 84.270 136.380 ;
        RECT 87.865 136.175 89.075 136.925 ;
        RECT 89.245 136.200 89.535 136.925 ;
        RECT 89.705 136.380 95.050 136.925 ;
        RECT 95.225 136.380 100.570 136.925 ;
        RECT 85.750 134.810 86.100 136.060 ;
        RECT 87.865 135.635 88.385 136.175 ;
        RECT 88.555 135.465 89.075 136.005 ;
        RECT 91.290 135.550 91.630 136.380 ;
        RECT 76.825 134.375 82.170 134.810 ;
        RECT 82.345 134.375 87.690 134.810 ;
        RECT 87.865 134.375 89.075 135.465 ;
        RECT 89.245 134.375 89.535 135.540 ;
        RECT 93.110 134.810 93.460 136.060 ;
        RECT 96.810 135.550 97.150 136.380 ;
        RECT 100.745 136.175 101.955 136.925 ;
        RECT 102.125 136.200 102.415 136.925 ;
        RECT 102.585 136.380 107.930 136.925 ;
        RECT 108.105 136.380 113.450 136.925 ;
        RECT 98.630 134.810 98.980 136.060 ;
        RECT 100.745 135.635 101.265 136.175 ;
        RECT 101.435 135.465 101.955 136.005 ;
        RECT 104.170 135.550 104.510 136.380 ;
        RECT 89.705 134.375 95.050 134.810 ;
        RECT 95.225 134.375 100.570 134.810 ;
        RECT 100.745 134.375 101.955 135.465 ;
        RECT 102.125 134.375 102.415 135.540 ;
        RECT 105.990 134.810 106.340 136.060 ;
        RECT 109.690 135.550 110.030 136.380 ;
        RECT 113.625 136.175 114.835 136.925 ;
        RECT 115.005 136.200 115.295 136.925 ;
        RECT 115.465 136.380 120.810 136.925 ;
        RECT 120.985 136.380 126.330 136.925 ;
        RECT 111.510 134.810 111.860 136.060 ;
        RECT 113.625 135.635 114.145 136.175 ;
        RECT 114.315 135.465 114.835 136.005 ;
        RECT 117.050 135.550 117.390 136.380 ;
        RECT 102.585 134.375 107.930 134.810 ;
        RECT 108.105 134.375 113.450 134.810 ;
        RECT 113.625 134.375 114.835 135.465 ;
        RECT 115.005 134.375 115.295 135.540 ;
        RECT 118.870 134.810 119.220 136.060 ;
        RECT 122.570 135.550 122.910 136.380 ;
        RECT 126.505 136.175 127.715 136.925 ;
        RECT 127.885 136.200 128.175 136.925 ;
        RECT 128.345 136.380 133.690 136.925 ;
        RECT 124.390 134.810 124.740 136.060 ;
        RECT 126.505 135.635 127.025 136.175 ;
        RECT 127.195 135.465 127.715 136.005 ;
        RECT 129.930 135.550 130.270 136.380 ;
        RECT 133.865 136.155 137.375 136.925 ;
        RECT 138.005 136.175 139.215 136.925 ;
        RECT 115.465 134.375 120.810 134.810 ;
        RECT 120.985 134.375 126.330 134.810 ;
        RECT 126.505 134.375 127.715 135.465 ;
        RECT 127.885 134.375 128.175 135.540 ;
        RECT 131.750 134.810 132.100 136.060 ;
        RECT 133.865 135.635 135.515 136.155 ;
        RECT 135.685 135.465 137.375 135.985 ;
        RECT 128.345 134.375 133.690 134.810 ;
        RECT 133.865 134.375 137.375 135.465 ;
        RECT 138.005 135.465 138.525 136.005 ;
        RECT 138.695 135.635 139.215 136.175 ;
        RECT 138.005 134.375 139.215 135.465 ;
        RECT 50.520 134.205 139.300 134.375 ;
        RECT 50.605 133.115 51.815 134.205 ;
        RECT 51.985 133.770 57.330 134.205 ;
        RECT 57.505 133.770 62.850 134.205 ;
        RECT 50.605 132.405 51.125 132.945 ;
        RECT 51.295 132.575 51.815 133.115 ;
        RECT 50.605 131.655 51.815 132.405 ;
        RECT 53.570 132.200 53.910 133.030 ;
        RECT 55.390 132.520 55.740 133.770 ;
        RECT 59.090 132.200 59.430 133.030 ;
        RECT 60.910 132.520 61.260 133.770 ;
        RECT 63.485 133.040 63.775 134.205 ;
        RECT 63.945 133.770 69.290 134.205 ;
        RECT 69.465 133.770 74.810 134.205 ;
        RECT 74.985 133.770 80.330 134.205 ;
        RECT 80.505 133.770 85.850 134.205 ;
        RECT 51.985 131.655 57.330 132.200 ;
        RECT 57.505 131.655 62.850 132.200 ;
        RECT 63.485 131.655 63.775 132.380 ;
        RECT 65.530 132.200 65.870 133.030 ;
        RECT 67.350 132.520 67.700 133.770 ;
        RECT 71.050 132.200 71.390 133.030 ;
        RECT 72.870 132.520 73.220 133.770 ;
        RECT 76.570 132.200 76.910 133.030 ;
        RECT 78.390 132.520 78.740 133.770 ;
        RECT 82.090 132.200 82.430 133.030 ;
        RECT 83.910 132.520 84.260 133.770 ;
        RECT 86.025 133.115 88.615 134.205 ;
        RECT 86.025 132.425 87.235 132.945 ;
        RECT 87.405 132.595 88.615 133.115 ;
        RECT 89.245 133.040 89.535 134.205 ;
        RECT 89.705 133.770 95.050 134.205 ;
        RECT 95.225 133.770 100.570 134.205 ;
        RECT 100.745 133.770 106.090 134.205 ;
        RECT 106.265 133.770 111.610 134.205 ;
        RECT 63.945 131.655 69.290 132.200 ;
        RECT 69.465 131.655 74.810 132.200 ;
        RECT 74.985 131.655 80.330 132.200 ;
        RECT 80.505 131.655 85.850 132.200 ;
        RECT 86.025 131.655 88.615 132.425 ;
        RECT 89.245 131.655 89.535 132.380 ;
        RECT 91.290 132.200 91.630 133.030 ;
        RECT 93.110 132.520 93.460 133.770 ;
        RECT 96.810 132.200 97.150 133.030 ;
        RECT 98.630 132.520 98.980 133.770 ;
        RECT 102.330 132.200 102.670 133.030 ;
        RECT 104.150 132.520 104.500 133.770 ;
        RECT 107.850 132.200 108.190 133.030 ;
        RECT 109.670 132.520 110.020 133.770 ;
        RECT 111.785 133.115 114.375 134.205 ;
        RECT 111.785 132.425 112.995 132.945 ;
        RECT 113.165 132.595 114.375 133.115 ;
        RECT 115.005 133.040 115.295 134.205 ;
        RECT 115.465 133.770 120.810 134.205 ;
        RECT 120.985 133.770 126.330 134.205 ;
        RECT 126.505 133.770 131.850 134.205 ;
        RECT 132.025 133.770 137.370 134.205 ;
        RECT 89.705 131.655 95.050 132.200 ;
        RECT 95.225 131.655 100.570 132.200 ;
        RECT 100.745 131.655 106.090 132.200 ;
        RECT 106.265 131.655 111.610 132.200 ;
        RECT 111.785 131.655 114.375 132.425 ;
        RECT 115.005 131.655 115.295 132.380 ;
        RECT 117.050 132.200 117.390 133.030 ;
        RECT 118.870 132.520 119.220 133.770 ;
        RECT 122.570 132.200 122.910 133.030 ;
        RECT 124.390 132.520 124.740 133.770 ;
        RECT 128.090 132.200 128.430 133.030 ;
        RECT 129.910 132.520 130.260 133.770 ;
        RECT 133.610 132.200 133.950 133.030 ;
        RECT 135.430 132.520 135.780 133.770 ;
        RECT 138.005 133.115 139.215 134.205 ;
        RECT 138.005 132.575 138.525 133.115 ;
        RECT 138.695 132.405 139.215 132.945 ;
        RECT 115.465 131.655 120.810 132.200 ;
        RECT 120.985 131.655 126.330 132.200 ;
        RECT 126.505 131.655 131.850 132.200 ;
        RECT 132.025 131.655 137.370 132.200 ;
        RECT 138.005 131.655 139.215 132.405 ;
        RECT 50.520 131.485 139.300 131.655 ;
        RECT 50.605 130.735 51.815 131.485 ;
        RECT 51.985 130.940 57.330 131.485 ;
        RECT 57.505 130.940 62.850 131.485 ;
        RECT 63.025 130.940 68.370 131.485 ;
        RECT 68.545 130.940 73.890 131.485 ;
        RECT 50.605 130.195 51.125 130.735 ;
        RECT 51.295 130.025 51.815 130.565 ;
        RECT 53.570 130.110 53.910 130.940 ;
        RECT 50.605 128.935 51.815 130.025 ;
        RECT 55.390 129.370 55.740 130.620 ;
        RECT 59.090 130.110 59.430 130.940 ;
        RECT 60.910 129.370 61.260 130.620 ;
        RECT 64.610 130.110 64.950 130.940 ;
        RECT 66.430 129.370 66.780 130.620 ;
        RECT 70.130 130.110 70.470 130.940 ;
        RECT 74.065 130.715 75.735 131.485 ;
        RECT 76.365 130.760 76.655 131.485 ;
        RECT 76.825 130.940 82.170 131.485 ;
        RECT 82.345 130.940 87.690 131.485 ;
        RECT 87.865 130.940 93.210 131.485 ;
        RECT 93.385 130.940 98.730 131.485 ;
        RECT 71.950 129.370 72.300 130.620 ;
        RECT 74.065 130.195 74.815 130.715 ;
        RECT 74.985 130.025 75.735 130.545 ;
        RECT 78.410 130.110 78.750 130.940 ;
        RECT 51.985 128.935 57.330 129.370 ;
        RECT 57.505 128.935 62.850 129.370 ;
        RECT 63.025 128.935 68.370 129.370 ;
        RECT 68.545 128.935 73.890 129.370 ;
        RECT 74.065 128.935 75.735 130.025 ;
        RECT 76.365 128.935 76.655 130.100 ;
        RECT 80.230 129.370 80.580 130.620 ;
        RECT 83.930 130.110 84.270 130.940 ;
        RECT 85.750 129.370 86.100 130.620 ;
        RECT 89.450 130.110 89.790 130.940 ;
        RECT 91.270 129.370 91.620 130.620 ;
        RECT 94.970 130.110 95.310 130.940 ;
        RECT 98.905 130.715 101.495 131.485 ;
        RECT 102.125 130.760 102.415 131.485 ;
        RECT 102.585 130.940 107.930 131.485 ;
        RECT 108.105 130.940 113.450 131.485 ;
        RECT 113.625 130.940 118.970 131.485 ;
        RECT 119.145 130.940 124.490 131.485 ;
        RECT 96.790 129.370 97.140 130.620 ;
        RECT 98.905 130.195 100.115 130.715 ;
        RECT 100.285 130.025 101.495 130.545 ;
        RECT 104.170 130.110 104.510 130.940 ;
        RECT 76.825 128.935 82.170 129.370 ;
        RECT 82.345 128.935 87.690 129.370 ;
        RECT 87.865 128.935 93.210 129.370 ;
        RECT 93.385 128.935 98.730 129.370 ;
        RECT 98.905 128.935 101.495 130.025 ;
        RECT 102.125 128.935 102.415 130.100 ;
        RECT 105.990 129.370 106.340 130.620 ;
        RECT 109.690 130.110 110.030 130.940 ;
        RECT 111.510 129.370 111.860 130.620 ;
        RECT 115.210 130.110 115.550 130.940 ;
        RECT 117.030 129.370 117.380 130.620 ;
        RECT 120.730 130.110 121.070 130.940 ;
        RECT 124.665 130.715 127.255 131.485 ;
        RECT 127.885 130.760 128.175 131.485 ;
        RECT 128.345 130.940 133.690 131.485 ;
        RECT 122.550 129.370 122.900 130.620 ;
        RECT 124.665 130.195 125.875 130.715 ;
        RECT 126.045 130.025 127.255 130.545 ;
        RECT 129.930 130.110 130.270 130.940 ;
        RECT 133.865 130.715 137.375 131.485 ;
        RECT 138.005 130.735 139.215 131.485 ;
        RECT 102.585 128.935 107.930 129.370 ;
        RECT 108.105 128.935 113.450 129.370 ;
        RECT 113.625 128.935 118.970 129.370 ;
        RECT 119.145 128.935 124.490 129.370 ;
        RECT 124.665 128.935 127.255 130.025 ;
        RECT 127.885 128.935 128.175 130.100 ;
        RECT 131.750 129.370 132.100 130.620 ;
        RECT 133.865 130.195 135.515 130.715 ;
        RECT 135.685 130.025 137.375 130.545 ;
        RECT 128.345 128.935 133.690 129.370 ;
        RECT 133.865 128.935 137.375 130.025 ;
        RECT 138.005 130.025 138.525 130.565 ;
        RECT 138.695 130.195 139.215 130.735 ;
        RECT 138.005 128.935 139.215 130.025 ;
        RECT 50.520 128.765 139.300 128.935 ;
        RECT 50.605 127.675 51.815 128.765 ;
        RECT 51.985 128.330 57.330 128.765 ;
        RECT 57.505 128.330 62.850 128.765 ;
        RECT 50.605 126.965 51.125 127.505 ;
        RECT 51.295 127.135 51.815 127.675 ;
        RECT 50.605 126.215 51.815 126.965 ;
        RECT 53.570 126.760 53.910 127.590 ;
        RECT 55.390 127.080 55.740 128.330 ;
        RECT 59.090 126.760 59.430 127.590 ;
        RECT 60.910 127.080 61.260 128.330 ;
        RECT 63.485 127.600 63.775 128.765 ;
        RECT 63.945 128.330 69.290 128.765 ;
        RECT 69.465 128.330 74.810 128.765 ;
        RECT 74.985 128.330 80.330 128.765 ;
        RECT 80.505 128.330 85.850 128.765 ;
        RECT 51.985 126.215 57.330 126.760 ;
        RECT 57.505 126.215 62.850 126.760 ;
        RECT 63.485 126.215 63.775 126.940 ;
        RECT 65.530 126.760 65.870 127.590 ;
        RECT 67.350 127.080 67.700 128.330 ;
        RECT 71.050 126.760 71.390 127.590 ;
        RECT 72.870 127.080 73.220 128.330 ;
        RECT 76.570 126.760 76.910 127.590 ;
        RECT 78.390 127.080 78.740 128.330 ;
        RECT 82.090 126.760 82.430 127.590 ;
        RECT 83.910 127.080 84.260 128.330 ;
        RECT 86.025 127.675 88.615 128.765 ;
        RECT 86.025 126.985 87.235 127.505 ;
        RECT 87.405 127.155 88.615 127.675 ;
        RECT 89.245 127.600 89.535 128.765 ;
        RECT 89.705 128.330 95.050 128.765 ;
        RECT 95.225 128.330 100.570 128.765 ;
        RECT 100.745 128.330 106.090 128.765 ;
        RECT 106.265 128.330 111.610 128.765 ;
        RECT 63.945 126.215 69.290 126.760 ;
        RECT 69.465 126.215 74.810 126.760 ;
        RECT 74.985 126.215 80.330 126.760 ;
        RECT 80.505 126.215 85.850 126.760 ;
        RECT 86.025 126.215 88.615 126.985 ;
        RECT 89.245 126.215 89.535 126.940 ;
        RECT 91.290 126.760 91.630 127.590 ;
        RECT 93.110 127.080 93.460 128.330 ;
        RECT 96.810 126.760 97.150 127.590 ;
        RECT 98.630 127.080 98.980 128.330 ;
        RECT 102.330 126.760 102.670 127.590 ;
        RECT 104.150 127.080 104.500 128.330 ;
        RECT 107.850 126.760 108.190 127.590 ;
        RECT 109.670 127.080 110.020 128.330 ;
        RECT 111.785 127.675 114.375 128.765 ;
        RECT 111.785 126.985 112.995 127.505 ;
        RECT 113.165 127.155 114.375 127.675 ;
        RECT 115.005 127.600 115.295 128.765 ;
        RECT 115.465 128.330 120.810 128.765 ;
        RECT 120.985 128.330 126.330 128.765 ;
        RECT 126.505 128.330 131.850 128.765 ;
        RECT 132.025 128.330 137.370 128.765 ;
        RECT 89.705 126.215 95.050 126.760 ;
        RECT 95.225 126.215 100.570 126.760 ;
        RECT 100.745 126.215 106.090 126.760 ;
        RECT 106.265 126.215 111.610 126.760 ;
        RECT 111.785 126.215 114.375 126.985 ;
        RECT 115.005 126.215 115.295 126.940 ;
        RECT 117.050 126.760 117.390 127.590 ;
        RECT 118.870 127.080 119.220 128.330 ;
        RECT 122.570 126.760 122.910 127.590 ;
        RECT 124.390 127.080 124.740 128.330 ;
        RECT 128.090 126.760 128.430 127.590 ;
        RECT 129.910 127.080 130.260 128.330 ;
        RECT 133.610 126.760 133.950 127.590 ;
        RECT 135.430 127.080 135.780 128.330 ;
        RECT 138.005 127.675 139.215 128.765 ;
        RECT 138.005 127.135 138.525 127.675 ;
        RECT 138.695 126.965 139.215 127.505 ;
        RECT 115.465 126.215 120.810 126.760 ;
        RECT 120.985 126.215 126.330 126.760 ;
        RECT 126.505 126.215 131.850 126.760 ;
        RECT 132.025 126.215 137.370 126.760 ;
        RECT 138.005 126.215 139.215 126.965 ;
        RECT 50.520 126.045 139.300 126.215 ;
        RECT 50.605 125.295 51.815 126.045 ;
        RECT 51.985 125.500 57.330 126.045 ;
        RECT 57.505 125.500 62.850 126.045 ;
        RECT 63.025 125.500 68.370 126.045 ;
        RECT 68.545 125.500 73.890 126.045 ;
        RECT 50.605 124.755 51.125 125.295 ;
        RECT 51.295 124.585 51.815 125.125 ;
        RECT 53.570 124.670 53.910 125.500 ;
        RECT 50.605 123.495 51.815 124.585 ;
        RECT 55.390 123.930 55.740 125.180 ;
        RECT 59.090 124.670 59.430 125.500 ;
        RECT 60.910 123.930 61.260 125.180 ;
        RECT 64.610 124.670 64.950 125.500 ;
        RECT 66.430 123.930 66.780 125.180 ;
        RECT 70.130 124.670 70.470 125.500 ;
        RECT 74.065 125.275 75.735 126.045 ;
        RECT 76.365 125.320 76.655 126.045 ;
        RECT 76.825 125.500 82.170 126.045 ;
        RECT 82.345 125.500 87.690 126.045 ;
        RECT 87.865 125.500 93.210 126.045 ;
        RECT 93.385 125.500 98.730 126.045 ;
        RECT 71.950 123.930 72.300 125.180 ;
        RECT 74.065 124.755 74.815 125.275 ;
        RECT 74.985 124.585 75.735 125.105 ;
        RECT 78.410 124.670 78.750 125.500 ;
        RECT 51.985 123.495 57.330 123.930 ;
        RECT 57.505 123.495 62.850 123.930 ;
        RECT 63.025 123.495 68.370 123.930 ;
        RECT 68.545 123.495 73.890 123.930 ;
        RECT 74.065 123.495 75.735 124.585 ;
        RECT 76.365 123.495 76.655 124.660 ;
        RECT 80.230 123.930 80.580 125.180 ;
        RECT 83.930 124.670 84.270 125.500 ;
        RECT 85.750 123.930 86.100 125.180 ;
        RECT 89.450 124.670 89.790 125.500 ;
        RECT 91.270 123.930 91.620 125.180 ;
        RECT 94.970 124.670 95.310 125.500 ;
        RECT 98.905 125.275 101.495 126.045 ;
        RECT 102.125 125.320 102.415 126.045 ;
        RECT 102.585 125.500 107.930 126.045 ;
        RECT 108.105 125.500 113.450 126.045 ;
        RECT 113.625 125.500 118.970 126.045 ;
        RECT 119.145 125.500 124.490 126.045 ;
        RECT 96.790 123.930 97.140 125.180 ;
        RECT 98.905 124.755 100.115 125.275 ;
        RECT 100.285 124.585 101.495 125.105 ;
        RECT 104.170 124.670 104.510 125.500 ;
        RECT 76.825 123.495 82.170 123.930 ;
        RECT 82.345 123.495 87.690 123.930 ;
        RECT 87.865 123.495 93.210 123.930 ;
        RECT 93.385 123.495 98.730 123.930 ;
        RECT 98.905 123.495 101.495 124.585 ;
        RECT 102.125 123.495 102.415 124.660 ;
        RECT 105.990 123.930 106.340 125.180 ;
        RECT 109.690 124.670 110.030 125.500 ;
        RECT 111.510 123.930 111.860 125.180 ;
        RECT 115.210 124.670 115.550 125.500 ;
        RECT 117.030 123.930 117.380 125.180 ;
        RECT 120.730 124.670 121.070 125.500 ;
        RECT 124.665 125.275 127.255 126.045 ;
        RECT 127.885 125.320 128.175 126.045 ;
        RECT 128.345 125.500 133.690 126.045 ;
        RECT 122.550 123.930 122.900 125.180 ;
        RECT 124.665 124.755 125.875 125.275 ;
        RECT 126.045 124.585 127.255 125.105 ;
        RECT 129.930 124.670 130.270 125.500 ;
        RECT 133.865 125.275 137.375 126.045 ;
        RECT 138.005 125.295 139.215 126.045 ;
        RECT 102.585 123.495 107.930 123.930 ;
        RECT 108.105 123.495 113.450 123.930 ;
        RECT 113.625 123.495 118.970 123.930 ;
        RECT 119.145 123.495 124.490 123.930 ;
        RECT 124.665 123.495 127.255 124.585 ;
        RECT 127.885 123.495 128.175 124.660 ;
        RECT 131.750 123.930 132.100 125.180 ;
        RECT 133.865 124.755 135.515 125.275 ;
        RECT 135.685 124.585 137.375 125.105 ;
        RECT 128.345 123.495 133.690 123.930 ;
        RECT 133.865 123.495 137.375 124.585 ;
        RECT 138.005 124.585 138.525 125.125 ;
        RECT 138.695 124.755 139.215 125.295 ;
        RECT 138.005 123.495 139.215 124.585 ;
        RECT 50.520 123.325 139.300 123.495 ;
        RECT 50.605 122.235 51.815 123.325 ;
        RECT 51.985 122.890 57.330 123.325 ;
        RECT 57.505 122.890 62.850 123.325 ;
        RECT 50.605 121.525 51.125 122.065 ;
        RECT 51.295 121.695 51.815 122.235 ;
        RECT 50.605 120.775 51.815 121.525 ;
        RECT 53.570 121.320 53.910 122.150 ;
        RECT 55.390 121.640 55.740 122.890 ;
        RECT 59.090 121.320 59.430 122.150 ;
        RECT 60.910 121.640 61.260 122.890 ;
        RECT 63.485 122.160 63.775 123.325 ;
        RECT 63.945 122.890 69.290 123.325 ;
        RECT 69.465 122.890 74.810 123.325 ;
        RECT 74.985 122.890 80.330 123.325 ;
        RECT 80.505 122.890 85.850 123.325 ;
        RECT 51.985 120.775 57.330 121.320 ;
        RECT 57.505 120.775 62.850 121.320 ;
        RECT 63.485 120.775 63.775 121.500 ;
        RECT 65.530 121.320 65.870 122.150 ;
        RECT 67.350 121.640 67.700 122.890 ;
        RECT 71.050 121.320 71.390 122.150 ;
        RECT 72.870 121.640 73.220 122.890 ;
        RECT 76.570 121.320 76.910 122.150 ;
        RECT 78.390 121.640 78.740 122.890 ;
        RECT 82.090 121.320 82.430 122.150 ;
        RECT 83.910 121.640 84.260 122.890 ;
        RECT 86.025 122.235 88.615 123.325 ;
        RECT 86.025 121.545 87.235 122.065 ;
        RECT 87.405 121.715 88.615 122.235 ;
        RECT 89.245 122.160 89.535 123.325 ;
        RECT 89.705 122.890 95.050 123.325 ;
        RECT 95.225 122.890 100.570 123.325 ;
        RECT 100.745 122.890 106.090 123.325 ;
        RECT 106.265 122.890 111.610 123.325 ;
        RECT 63.945 120.775 69.290 121.320 ;
        RECT 69.465 120.775 74.810 121.320 ;
        RECT 74.985 120.775 80.330 121.320 ;
        RECT 80.505 120.775 85.850 121.320 ;
        RECT 86.025 120.775 88.615 121.545 ;
        RECT 89.245 120.775 89.535 121.500 ;
        RECT 91.290 121.320 91.630 122.150 ;
        RECT 93.110 121.640 93.460 122.890 ;
        RECT 96.810 121.320 97.150 122.150 ;
        RECT 98.630 121.640 98.980 122.890 ;
        RECT 102.330 121.320 102.670 122.150 ;
        RECT 104.150 121.640 104.500 122.890 ;
        RECT 107.850 121.320 108.190 122.150 ;
        RECT 109.670 121.640 110.020 122.890 ;
        RECT 111.785 122.235 114.375 123.325 ;
        RECT 111.785 121.545 112.995 122.065 ;
        RECT 113.165 121.715 114.375 122.235 ;
        RECT 115.005 122.160 115.295 123.325 ;
        RECT 115.465 122.890 120.810 123.325 ;
        RECT 120.985 122.890 126.330 123.325 ;
        RECT 126.505 122.890 131.850 123.325 ;
        RECT 132.025 122.890 137.370 123.325 ;
        RECT 89.705 120.775 95.050 121.320 ;
        RECT 95.225 120.775 100.570 121.320 ;
        RECT 100.745 120.775 106.090 121.320 ;
        RECT 106.265 120.775 111.610 121.320 ;
        RECT 111.785 120.775 114.375 121.545 ;
        RECT 115.005 120.775 115.295 121.500 ;
        RECT 117.050 121.320 117.390 122.150 ;
        RECT 118.870 121.640 119.220 122.890 ;
        RECT 122.570 121.320 122.910 122.150 ;
        RECT 124.390 121.640 124.740 122.890 ;
        RECT 128.090 121.320 128.430 122.150 ;
        RECT 129.910 121.640 130.260 122.890 ;
        RECT 133.610 121.320 133.950 122.150 ;
        RECT 135.430 121.640 135.780 122.890 ;
        RECT 138.005 122.235 139.215 123.325 ;
        RECT 138.005 121.695 138.525 122.235 ;
        RECT 138.695 121.525 139.215 122.065 ;
        RECT 115.465 120.775 120.810 121.320 ;
        RECT 120.985 120.775 126.330 121.320 ;
        RECT 126.505 120.775 131.850 121.320 ;
        RECT 132.025 120.775 137.370 121.320 ;
        RECT 138.005 120.775 139.215 121.525 ;
        RECT 50.520 120.605 139.300 120.775 ;
        RECT 50.605 119.855 51.815 120.605 ;
        RECT 51.985 120.060 57.330 120.605 ;
        RECT 57.505 120.060 62.850 120.605 ;
        RECT 63.025 120.060 68.370 120.605 ;
        RECT 68.545 120.060 73.890 120.605 ;
        RECT 50.605 119.315 51.125 119.855 ;
        RECT 51.295 119.145 51.815 119.685 ;
        RECT 53.570 119.230 53.910 120.060 ;
        RECT 50.605 118.055 51.815 119.145 ;
        RECT 55.390 118.490 55.740 119.740 ;
        RECT 59.090 119.230 59.430 120.060 ;
        RECT 60.910 118.490 61.260 119.740 ;
        RECT 64.610 119.230 64.950 120.060 ;
        RECT 66.430 118.490 66.780 119.740 ;
        RECT 70.130 119.230 70.470 120.060 ;
        RECT 74.065 119.835 75.735 120.605 ;
        RECT 76.365 119.880 76.655 120.605 ;
        RECT 76.825 120.060 82.170 120.605 ;
        RECT 82.345 120.060 87.690 120.605 ;
        RECT 87.865 120.060 93.210 120.605 ;
        RECT 93.385 120.060 98.730 120.605 ;
        RECT 71.950 118.490 72.300 119.740 ;
        RECT 74.065 119.315 74.815 119.835 ;
        RECT 74.985 119.145 75.735 119.665 ;
        RECT 78.410 119.230 78.750 120.060 ;
        RECT 51.985 118.055 57.330 118.490 ;
        RECT 57.505 118.055 62.850 118.490 ;
        RECT 63.025 118.055 68.370 118.490 ;
        RECT 68.545 118.055 73.890 118.490 ;
        RECT 74.065 118.055 75.735 119.145 ;
        RECT 76.365 118.055 76.655 119.220 ;
        RECT 80.230 118.490 80.580 119.740 ;
        RECT 83.930 119.230 84.270 120.060 ;
        RECT 85.750 118.490 86.100 119.740 ;
        RECT 89.450 119.230 89.790 120.060 ;
        RECT 91.270 118.490 91.620 119.740 ;
        RECT 94.970 119.230 95.310 120.060 ;
        RECT 98.905 119.835 101.495 120.605 ;
        RECT 102.125 119.880 102.415 120.605 ;
        RECT 102.585 120.060 107.930 120.605 ;
        RECT 108.105 120.060 113.450 120.605 ;
        RECT 113.625 120.060 118.970 120.605 ;
        RECT 119.145 120.060 124.490 120.605 ;
        RECT 96.790 118.490 97.140 119.740 ;
        RECT 98.905 119.315 100.115 119.835 ;
        RECT 100.285 119.145 101.495 119.665 ;
        RECT 104.170 119.230 104.510 120.060 ;
        RECT 76.825 118.055 82.170 118.490 ;
        RECT 82.345 118.055 87.690 118.490 ;
        RECT 87.865 118.055 93.210 118.490 ;
        RECT 93.385 118.055 98.730 118.490 ;
        RECT 98.905 118.055 101.495 119.145 ;
        RECT 102.125 118.055 102.415 119.220 ;
        RECT 105.990 118.490 106.340 119.740 ;
        RECT 109.690 119.230 110.030 120.060 ;
        RECT 111.510 118.490 111.860 119.740 ;
        RECT 115.210 119.230 115.550 120.060 ;
        RECT 117.030 118.490 117.380 119.740 ;
        RECT 120.730 119.230 121.070 120.060 ;
        RECT 124.665 119.835 127.255 120.605 ;
        RECT 127.885 119.880 128.175 120.605 ;
        RECT 128.345 120.060 133.690 120.605 ;
        RECT 122.550 118.490 122.900 119.740 ;
        RECT 124.665 119.315 125.875 119.835 ;
        RECT 126.045 119.145 127.255 119.665 ;
        RECT 129.930 119.230 130.270 120.060 ;
        RECT 133.865 119.835 137.375 120.605 ;
        RECT 138.005 119.855 139.215 120.605 ;
        RECT 102.585 118.055 107.930 118.490 ;
        RECT 108.105 118.055 113.450 118.490 ;
        RECT 113.625 118.055 118.970 118.490 ;
        RECT 119.145 118.055 124.490 118.490 ;
        RECT 124.665 118.055 127.255 119.145 ;
        RECT 127.885 118.055 128.175 119.220 ;
        RECT 131.750 118.490 132.100 119.740 ;
        RECT 133.865 119.315 135.515 119.835 ;
        RECT 135.685 119.145 137.375 119.665 ;
        RECT 128.345 118.055 133.690 118.490 ;
        RECT 133.865 118.055 137.375 119.145 ;
        RECT 138.005 119.145 138.525 119.685 ;
        RECT 138.695 119.315 139.215 119.855 ;
        RECT 138.005 118.055 139.215 119.145 ;
        RECT 50.520 117.885 139.300 118.055 ;
        RECT 50.605 116.795 51.815 117.885 ;
        RECT 51.985 117.450 57.330 117.885 ;
        RECT 57.505 117.450 62.850 117.885 ;
        RECT 50.605 116.085 51.125 116.625 ;
        RECT 51.295 116.255 51.815 116.795 ;
        RECT 50.605 115.335 51.815 116.085 ;
        RECT 53.570 115.880 53.910 116.710 ;
        RECT 55.390 116.200 55.740 117.450 ;
        RECT 59.090 115.880 59.430 116.710 ;
        RECT 60.910 116.200 61.260 117.450 ;
        RECT 63.485 116.720 63.775 117.885 ;
        RECT 63.945 117.450 69.290 117.885 ;
        RECT 69.465 117.450 74.810 117.885 ;
        RECT 74.985 117.450 80.330 117.885 ;
        RECT 80.505 117.450 85.850 117.885 ;
        RECT 51.985 115.335 57.330 115.880 ;
        RECT 57.505 115.335 62.850 115.880 ;
        RECT 63.485 115.335 63.775 116.060 ;
        RECT 65.530 115.880 65.870 116.710 ;
        RECT 67.350 116.200 67.700 117.450 ;
        RECT 71.050 115.880 71.390 116.710 ;
        RECT 72.870 116.200 73.220 117.450 ;
        RECT 76.570 115.880 76.910 116.710 ;
        RECT 78.390 116.200 78.740 117.450 ;
        RECT 82.090 115.880 82.430 116.710 ;
        RECT 83.910 116.200 84.260 117.450 ;
        RECT 86.025 116.795 88.615 117.885 ;
        RECT 86.025 116.105 87.235 116.625 ;
        RECT 87.405 116.275 88.615 116.795 ;
        RECT 89.245 116.720 89.535 117.885 ;
        RECT 89.705 117.450 95.050 117.885 ;
        RECT 95.225 117.450 100.570 117.885 ;
        RECT 100.745 117.450 106.090 117.885 ;
        RECT 106.265 117.450 111.610 117.885 ;
        RECT 63.945 115.335 69.290 115.880 ;
        RECT 69.465 115.335 74.810 115.880 ;
        RECT 74.985 115.335 80.330 115.880 ;
        RECT 80.505 115.335 85.850 115.880 ;
        RECT 86.025 115.335 88.615 116.105 ;
        RECT 89.245 115.335 89.535 116.060 ;
        RECT 91.290 115.880 91.630 116.710 ;
        RECT 93.110 116.200 93.460 117.450 ;
        RECT 96.810 115.880 97.150 116.710 ;
        RECT 98.630 116.200 98.980 117.450 ;
        RECT 102.330 115.880 102.670 116.710 ;
        RECT 104.150 116.200 104.500 117.450 ;
        RECT 107.850 115.880 108.190 116.710 ;
        RECT 109.670 116.200 110.020 117.450 ;
        RECT 111.785 116.795 114.375 117.885 ;
        RECT 111.785 116.105 112.995 116.625 ;
        RECT 113.165 116.275 114.375 116.795 ;
        RECT 115.005 116.720 115.295 117.885 ;
        RECT 115.465 117.450 120.810 117.885 ;
        RECT 120.985 117.450 126.330 117.885 ;
        RECT 126.505 117.450 131.850 117.885 ;
        RECT 132.025 117.450 137.370 117.885 ;
        RECT 89.705 115.335 95.050 115.880 ;
        RECT 95.225 115.335 100.570 115.880 ;
        RECT 100.745 115.335 106.090 115.880 ;
        RECT 106.265 115.335 111.610 115.880 ;
        RECT 111.785 115.335 114.375 116.105 ;
        RECT 115.005 115.335 115.295 116.060 ;
        RECT 117.050 115.880 117.390 116.710 ;
        RECT 118.870 116.200 119.220 117.450 ;
        RECT 122.570 115.880 122.910 116.710 ;
        RECT 124.390 116.200 124.740 117.450 ;
        RECT 128.090 115.880 128.430 116.710 ;
        RECT 129.910 116.200 130.260 117.450 ;
        RECT 133.610 115.880 133.950 116.710 ;
        RECT 135.430 116.200 135.780 117.450 ;
        RECT 138.005 116.795 139.215 117.885 ;
        RECT 138.005 116.255 138.525 116.795 ;
        RECT 138.695 116.085 139.215 116.625 ;
        RECT 115.465 115.335 120.810 115.880 ;
        RECT 120.985 115.335 126.330 115.880 ;
        RECT 126.505 115.335 131.850 115.880 ;
        RECT 132.025 115.335 137.370 115.880 ;
        RECT 138.005 115.335 139.215 116.085 ;
        RECT 50.520 115.165 139.300 115.335 ;
        RECT 50.605 114.415 51.815 115.165 ;
        RECT 51.985 114.620 57.330 115.165 ;
        RECT 57.505 114.620 62.850 115.165 ;
        RECT 63.025 114.620 68.370 115.165 ;
        RECT 68.545 114.620 73.890 115.165 ;
        RECT 50.605 113.875 51.125 114.415 ;
        RECT 51.295 113.705 51.815 114.245 ;
        RECT 53.570 113.790 53.910 114.620 ;
        RECT 50.605 112.615 51.815 113.705 ;
        RECT 55.390 113.050 55.740 114.300 ;
        RECT 59.090 113.790 59.430 114.620 ;
        RECT 60.910 113.050 61.260 114.300 ;
        RECT 64.610 113.790 64.950 114.620 ;
        RECT 66.430 113.050 66.780 114.300 ;
        RECT 70.130 113.790 70.470 114.620 ;
        RECT 74.065 114.395 75.735 115.165 ;
        RECT 76.365 114.440 76.655 115.165 ;
        RECT 76.825 114.620 82.170 115.165 ;
        RECT 82.345 114.620 87.690 115.165 ;
        RECT 87.865 114.620 93.210 115.165 ;
        RECT 93.385 114.620 98.730 115.165 ;
        RECT 71.950 113.050 72.300 114.300 ;
        RECT 74.065 113.875 74.815 114.395 ;
        RECT 74.985 113.705 75.735 114.225 ;
        RECT 78.410 113.790 78.750 114.620 ;
        RECT 51.985 112.615 57.330 113.050 ;
        RECT 57.505 112.615 62.850 113.050 ;
        RECT 63.025 112.615 68.370 113.050 ;
        RECT 68.545 112.615 73.890 113.050 ;
        RECT 74.065 112.615 75.735 113.705 ;
        RECT 76.365 112.615 76.655 113.780 ;
        RECT 80.230 113.050 80.580 114.300 ;
        RECT 83.930 113.790 84.270 114.620 ;
        RECT 85.750 113.050 86.100 114.300 ;
        RECT 89.450 113.790 89.790 114.620 ;
        RECT 91.270 113.050 91.620 114.300 ;
        RECT 94.970 113.790 95.310 114.620 ;
        RECT 98.905 114.395 101.495 115.165 ;
        RECT 102.125 114.440 102.415 115.165 ;
        RECT 102.585 114.620 107.930 115.165 ;
        RECT 108.105 114.620 113.450 115.165 ;
        RECT 113.625 114.620 118.970 115.165 ;
        RECT 119.145 114.620 124.490 115.165 ;
        RECT 96.790 113.050 97.140 114.300 ;
        RECT 98.905 113.875 100.115 114.395 ;
        RECT 100.285 113.705 101.495 114.225 ;
        RECT 104.170 113.790 104.510 114.620 ;
        RECT 76.825 112.615 82.170 113.050 ;
        RECT 82.345 112.615 87.690 113.050 ;
        RECT 87.865 112.615 93.210 113.050 ;
        RECT 93.385 112.615 98.730 113.050 ;
        RECT 98.905 112.615 101.495 113.705 ;
        RECT 102.125 112.615 102.415 113.780 ;
        RECT 105.990 113.050 106.340 114.300 ;
        RECT 109.690 113.790 110.030 114.620 ;
        RECT 111.510 113.050 111.860 114.300 ;
        RECT 115.210 113.790 115.550 114.620 ;
        RECT 117.030 113.050 117.380 114.300 ;
        RECT 120.730 113.790 121.070 114.620 ;
        RECT 124.665 114.395 127.255 115.165 ;
        RECT 127.885 114.440 128.175 115.165 ;
        RECT 128.345 114.620 133.690 115.165 ;
        RECT 122.550 113.050 122.900 114.300 ;
        RECT 124.665 113.875 125.875 114.395 ;
        RECT 126.045 113.705 127.255 114.225 ;
        RECT 129.930 113.790 130.270 114.620 ;
        RECT 133.865 114.395 137.375 115.165 ;
        RECT 138.005 114.415 139.215 115.165 ;
        RECT 102.585 112.615 107.930 113.050 ;
        RECT 108.105 112.615 113.450 113.050 ;
        RECT 113.625 112.615 118.970 113.050 ;
        RECT 119.145 112.615 124.490 113.050 ;
        RECT 124.665 112.615 127.255 113.705 ;
        RECT 127.885 112.615 128.175 113.780 ;
        RECT 131.750 113.050 132.100 114.300 ;
        RECT 133.865 113.875 135.515 114.395 ;
        RECT 135.685 113.705 137.375 114.225 ;
        RECT 128.345 112.615 133.690 113.050 ;
        RECT 133.865 112.615 137.375 113.705 ;
        RECT 138.005 113.705 138.525 114.245 ;
        RECT 138.695 113.875 139.215 114.415 ;
        RECT 138.005 112.615 139.215 113.705 ;
        RECT 50.520 112.445 139.300 112.615 ;
        RECT 50.605 111.355 51.815 112.445 ;
        RECT 51.985 112.010 57.330 112.445 ;
        RECT 57.505 112.010 62.850 112.445 ;
        RECT 50.605 110.645 51.125 111.185 ;
        RECT 51.295 110.815 51.815 111.355 ;
        RECT 50.605 109.895 51.815 110.645 ;
        RECT 53.570 110.440 53.910 111.270 ;
        RECT 55.390 110.760 55.740 112.010 ;
        RECT 59.090 110.440 59.430 111.270 ;
        RECT 60.910 110.760 61.260 112.010 ;
        RECT 63.485 111.280 63.775 112.445 ;
        RECT 63.945 112.010 69.290 112.445 ;
        RECT 69.465 112.010 74.810 112.445 ;
        RECT 74.985 112.010 80.330 112.445 ;
        RECT 80.505 112.010 85.850 112.445 ;
        RECT 51.985 109.895 57.330 110.440 ;
        RECT 57.505 109.895 62.850 110.440 ;
        RECT 63.485 109.895 63.775 110.620 ;
        RECT 65.530 110.440 65.870 111.270 ;
        RECT 67.350 110.760 67.700 112.010 ;
        RECT 71.050 110.440 71.390 111.270 ;
        RECT 72.870 110.760 73.220 112.010 ;
        RECT 76.570 110.440 76.910 111.270 ;
        RECT 78.390 110.760 78.740 112.010 ;
        RECT 82.090 110.440 82.430 111.270 ;
        RECT 83.910 110.760 84.260 112.010 ;
        RECT 86.025 111.355 88.615 112.445 ;
        RECT 86.025 110.665 87.235 111.185 ;
        RECT 87.405 110.835 88.615 111.355 ;
        RECT 89.245 111.280 89.535 112.445 ;
        RECT 89.705 112.010 95.050 112.445 ;
        RECT 95.225 112.010 100.570 112.445 ;
        RECT 100.745 112.010 106.090 112.445 ;
        RECT 106.265 112.010 111.610 112.445 ;
        RECT 63.945 109.895 69.290 110.440 ;
        RECT 69.465 109.895 74.810 110.440 ;
        RECT 74.985 109.895 80.330 110.440 ;
        RECT 80.505 109.895 85.850 110.440 ;
        RECT 86.025 109.895 88.615 110.665 ;
        RECT 89.245 109.895 89.535 110.620 ;
        RECT 91.290 110.440 91.630 111.270 ;
        RECT 93.110 110.760 93.460 112.010 ;
        RECT 96.810 110.440 97.150 111.270 ;
        RECT 98.630 110.760 98.980 112.010 ;
        RECT 102.330 110.440 102.670 111.270 ;
        RECT 104.150 110.760 104.500 112.010 ;
        RECT 107.850 110.440 108.190 111.270 ;
        RECT 109.670 110.760 110.020 112.010 ;
        RECT 111.785 111.355 114.375 112.445 ;
        RECT 111.785 110.665 112.995 111.185 ;
        RECT 113.165 110.835 114.375 111.355 ;
        RECT 115.005 111.280 115.295 112.445 ;
        RECT 115.465 112.010 120.810 112.445 ;
        RECT 120.985 112.010 126.330 112.445 ;
        RECT 126.505 112.010 131.850 112.445 ;
        RECT 132.025 112.010 137.370 112.445 ;
        RECT 89.705 109.895 95.050 110.440 ;
        RECT 95.225 109.895 100.570 110.440 ;
        RECT 100.745 109.895 106.090 110.440 ;
        RECT 106.265 109.895 111.610 110.440 ;
        RECT 111.785 109.895 114.375 110.665 ;
        RECT 115.005 109.895 115.295 110.620 ;
        RECT 117.050 110.440 117.390 111.270 ;
        RECT 118.870 110.760 119.220 112.010 ;
        RECT 122.570 110.440 122.910 111.270 ;
        RECT 124.390 110.760 124.740 112.010 ;
        RECT 128.090 110.440 128.430 111.270 ;
        RECT 129.910 110.760 130.260 112.010 ;
        RECT 133.610 110.440 133.950 111.270 ;
        RECT 135.430 110.760 135.780 112.010 ;
        RECT 138.005 111.355 139.215 112.445 ;
        RECT 138.005 110.815 138.525 111.355 ;
        RECT 138.695 110.645 139.215 111.185 ;
        RECT 115.465 109.895 120.810 110.440 ;
        RECT 120.985 109.895 126.330 110.440 ;
        RECT 126.505 109.895 131.850 110.440 ;
        RECT 132.025 109.895 137.370 110.440 ;
        RECT 138.005 109.895 139.215 110.645 ;
        RECT 50.520 109.725 139.300 109.895 ;
        RECT 50.605 108.975 51.815 109.725 ;
        RECT 51.985 109.180 57.330 109.725 ;
        RECT 57.505 109.180 62.850 109.725 ;
        RECT 50.605 108.435 51.125 108.975 ;
        RECT 51.295 108.265 51.815 108.805 ;
        RECT 53.570 108.350 53.910 109.180 ;
        RECT 50.605 107.175 51.815 108.265 ;
        RECT 55.390 107.610 55.740 108.860 ;
        RECT 59.090 108.350 59.430 109.180 ;
        RECT 63.025 108.955 64.695 109.725 ;
        RECT 60.910 107.610 61.260 108.860 ;
        RECT 63.025 108.435 63.775 108.955 ;
        RECT 65.365 108.905 65.595 109.725 ;
        RECT 65.765 108.925 66.095 109.555 ;
        RECT 63.945 108.265 64.695 108.785 ;
        RECT 65.345 108.485 65.675 108.735 ;
        RECT 65.845 108.325 66.095 108.925 ;
        RECT 66.265 108.905 66.475 109.725 ;
        RECT 66.795 109.175 66.965 109.555 ;
        RECT 67.180 109.345 67.510 109.725 ;
        RECT 66.795 109.005 67.510 109.175 ;
        RECT 66.705 108.455 67.060 108.825 ;
        RECT 67.340 108.815 67.510 109.005 ;
        RECT 67.680 108.980 67.935 109.555 ;
        RECT 67.340 108.485 67.595 108.815 ;
        RECT 51.985 107.175 57.330 107.610 ;
        RECT 57.505 107.175 62.850 107.610 ;
        RECT 63.025 107.175 64.695 108.265 ;
        RECT 65.365 107.175 65.595 108.315 ;
        RECT 65.765 107.345 66.095 108.325 ;
        RECT 66.265 107.175 66.475 108.315 ;
        RECT 67.340 108.275 67.510 108.485 ;
        RECT 66.795 108.105 67.510 108.275 ;
        RECT 67.765 108.250 67.935 108.980 ;
        RECT 68.110 108.885 68.370 109.725 ;
        RECT 68.545 109.180 73.890 109.725 ;
        RECT 70.130 108.350 70.470 109.180 ;
        RECT 74.065 108.955 75.735 109.725 ;
        RECT 76.365 109.000 76.655 109.725 ;
        RECT 76.825 109.180 82.170 109.725 ;
        RECT 82.345 109.180 87.690 109.725 ;
        RECT 87.865 109.180 93.210 109.725 ;
        RECT 93.385 109.180 98.730 109.725 ;
        RECT 66.795 107.345 66.965 108.105 ;
        RECT 67.180 107.175 67.510 107.935 ;
        RECT 67.680 107.345 67.935 108.250 ;
        RECT 68.110 107.175 68.370 108.325 ;
        RECT 71.950 107.610 72.300 108.860 ;
        RECT 74.065 108.435 74.815 108.955 ;
        RECT 74.985 108.265 75.735 108.785 ;
        RECT 78.410 108.350 78.750 109.180 ;
        RECT 68.545 107.175 73.890 107.610 ;
        RECT 74.065 107.175 75.735 108.265 ;
        RECT 76.365 107.175 76.655 108.340 ;
        RECT 80.230 107.610 80.580 108.860 ;
        RECT 83.930 108.350 84.270 109.180 ;
        RECT 85.750 107.610 86.100 108.860 ;
        RECT 89.450 108.350 89.790 109.180 ;
        RECT 91.270 107.610 91.620 108.860 ;
        RECT 94.970 108.350 95.310 109.180 ;
        RECT 98.905 108.955 101.495 109.725 ;
        RECT 102.125 109.000 102.415 109.725 ;
        RECT 102.585 109.180 107.930 109.725 ;
        RECT 108.105 109.180 113.450 109.725 ;
        RECT 113.625 109.180 118.970 109.725 ;
        RECT 119.145 109.180 124.490 109.725 ;
        RECT 96.790 107.610 97.140 108.860 ;
        RECT 98.905 108.435 100.115 108.955 ;
        RECT 100.285 108.265 101.495 108.785 ;
        RECT 104.170 108.350 104.510 109.180 ;
        RECT 76.825 107.175 82.170 107.610 ;
        RECT 82.345 107.175 87.690 107.610 ;
        RECT 87.865 107.175 93.210 107.610 ;
        RECT 93.385 107.175 98.730 107.610 ;
        RECT 98.905 107.175 101.495 108.265 ;
        RECT 102.125 107.175 102.415 108.340 ;
        RECT 105.990 107.610 106.340 108.860 ;
        RECT 109.690 108.350 110.030 109.180 ;
        RECT 111.510 107.610 111.860 108.860 ;
        RECT 115.210 108.350 115.550 109.180 ;
        RECT 117.030 107.610 117.380 108.860 ;
        RECT 120.730 108.350 121.070 109.180 ;
        RECT 124.665 108.955 127.255 109.725 ;
        RECT 127.885 109.000 128.175 109.725 ;
        RECT 128.345 109.180 133.690 109.725 ;
        RECT 122.550 107.610 122.900 108.860 ;
        RECT 124.665 108.435 125.875 108.955 ;
        RECT 126.045 108.265 127.255 108.785 ;
        RECT 129.930 108.350 130.270 109.180 ;
        RECT 133.865 108.955 137.375 109.725 ;
        RECT 138.005 108.975 139.215 109.725 ;
        RECT 102.585 107.175 107.930 107.610 ;
        RECT 108.105 107.175 113.450 107.610 ;
        RECT 113.625 107.175 118.970 107.610 ;
        RECT 119.145 107.175 124.490 107.610 ;
        RECT 124.665 107.175 127.255 108.265 ;
        RECT 127.885 107.175 128.175 108.340 ;
        RECT 131.750 107.610 132.100 108.860 ;
        RECT 133.865 108.435 135.515 108.955 ;
        RECT 135.685 108.265 137.375 108.785 ;
        RECT 128.345 107.175 133.690 107.610 ;
        RECT 133.865 107.175 137.375 108.265 ;
        RECT 138.005 108.265 138.525 108.805 ;
        RECT 138.695 108.435 139.215 108.975 ;
        RECT 138.005 107.175 139.215 108.265 ;
        RECT 50.520 107.005 139.300 107.175 ;
        RECT 50.605 105.915 51.815 107.005 ;
        RECT 51.985 105.915 55.495 107.005 ;
        RECT 50.605 105.205 51.125 105.745 ;
        RECT 51.295 105.375 51.815 105.915 ;
        RECT 51.985 105.225 53.635 105.745 ;
        RECT 53.805 105.395 55.495 105.915 ;
        RECT 56.185 105.865 56.395 107.005 ;
        RECT 56.565 105.855 56.895 106.835 ;
        RECT 57.065 105.865 57.295 107.005 ;
        RECT 57.505 105.865 57.785 107.005 ;
        RECT 57.955 105.855 58.285 106.835 ;
        RECT 58.455 105.865 58.715 107.005 ;
        RECT 58.885 105.865 60.505 106.835 ;
        RECT 60.675 106.545 61.040 107.005 ;
        RECT 61.210 106.375 61.465 106.830 ;
        RECT 61.635 106.545 61.965 107.005 ;
        RECT 62.135 106.375 62.395 106.835 ;
        RECT 60.675 106.170 61.465 106.375 ;
        RECT 50.605 104.455 51.815 105.205 ;
        RECT 51.985 104.455 55.495 105.225 ;
        RECT 56.185 104.455 56.395 105.275 ;
        RECT 56.565 105.255 56.815 105.855 ;
        RECT 58.020 105.815 58.195 105.855 ;
        RECT 56.985 105.445 57.315 105.695 ;
        RECT 57.515 105.425 57.850 105.695 ;
        RECT 56.565 104.625 56.895 105.255 ;
        RECT 57.065 104.455 57.295 105.275 ;
        RECT 58.020 105.255 58.190 105.815 ;
        RECT 58.360 105.445 58.695 105.695 ;
        RECT 57.505 104.455 57.815 105.255 ;
        RECT 58.020 104.625 58.715 105.255 ;
        RECT 58.885 105.195 59.225 105.865 ;
        RECT 60.675 105.695 61.070 106.170 ;
        RECT 61.740 106.155 62.395 106.375 ;
        RECT 59.395 105.365 59.775 105.695 ;
        RECT 59.945 105.445 61.070 105.695 ;
        RECT 61.240 105.445 61.570 106.000 ;
        RECT 59.525 105.275 59.775 105.365 ;
        RECT 58.885 104.625 59.355 105.195 ;
        RECT 59.525 105.105 60.625 105.275 ;
        RECT 59.525 104.455 60.285 104.935 ;
        RECT 60.455 104.835 60.625 105.105 ;
        RECT 60.795 105.255 61.070 105.445 ;
        RECT 60.795 105.005 61.125 105.255 ;
        RECT 61.740 105.195 61.955 106.155 ;
        RECT 62.125 105.365 62.395 105.985 ;
        RECT 63.485 105.840 63.775 107.005 ;
        RECT 63.945 106.570 69.290 107.005 ;
        RECT 69.465 106.570 74.810 107.005 ;
        RECT 74.985 106.570 80.330 107.005 ;
        RECT 80.505 106.570 85.850 107.005 ;
        RECT 61.295 104.985 62.395 105.195 ;
        RECT 61.295 104.835 61.465 104.985 ;
        RECT 60.455 104.625 61.465 104.835 ;
        RECT 61.635 104.455 61.965 104.815 ;
        RECT 62.135 104.650 62.395 104.985 ;
        RECT 63.485 104.455 63.775 105.180 ;
        RECT 65.530 105.000 65.870 105.830 ;
        RECT 67.350 105.320 67.700 106.570 ;
        RECT 71.050 105.000 71.390 105.830 ;
        RECT 72.870 105.320 73.220 106.570 ;
        RECT 76.570 105.000 76.910 105.830 ;
        RECT 78.390 105.320 78.740 106.570 ;
        RECT 82.090 105.000 82.430 105.830 ;
        RECT 83.910 105.320 84.260 106.570 ;
        RECT 86.025 105.915 88.615 107.005 ;
        RECT 86.025 105.225 87.235 105.745 ;
        RECT 87.405 105.395 88.615 105.915 ;
        RECT 89.245 105.840 89.535 107.005 ;
        RECT 89.705 106.570 95.050 107.005 ;
        RECT 95.225 106.570 100.570 107.005 ;
        RECT 100.745 106.570 106.090 107.005 ;
        RECT 106.265 106.570 111.610 107.005 ;
        RECT 63.945 104.455 69.290 105.000 ;
        RECT 69.465 104.455 74.810 105.000 ;
        RECT 74.985 104.455 80.330 105.000 ;
        RECT 80.505 104.455 85.850 105.000 ;
        RECT 86.025 104.455 88.615 105.225 ;
        RECT 89.245 104.455 89.535 105.180 ;
        RECT 91.290 105.000 91.630 105.830 ;
        RECT 93.110 105.320 93.460 106.570 ;
        RECT 96.810 105.000 97.150 105.830 ;
        RECT 98.630 105.320 98.980 106.570 ;
        RECT 102.330 105.000 102.670 105.830 ;
        RECT 104.150 105.320 104.500 106.570 ;
        RECT 107.850 105.000 108.190 105.830 ;
        RECT 109.670 105.320 110.020 106.570 ;
        RECT 111.785 105.915 114.375 107.005 ;
        RECT 111.785 105.225 112.995 105.745 ;
        RECT 113.165 105.395 114.375 105.915 ;
        RECT 115.005 105.840 115.295 107.005 ;
        RECT 115.465 106.570 120.810 107.005 ;
        RECT 120.985 106.570 126.330 107.005 ;
        RECT 126.505 106.570 131.850 107.005 ;
        RECT 132.025 106.570 137.370 107.005 ;
        RECT 89.705 104.455 95.050 105.000 ;
        RECT 95.225 104.455 100.570 105.000 ;
        RECT 100.745 104.455 106.090 105.000 ;
        RECT 106.265 104.455 111.610 105.000 ;
        RECT 111.785 104.455 114.375 105.225 ;
        RECT 115.005 104.455 115.295 105.180 ;
        RECT 117.050 105.000 117.390 105.830 ;
        RECT 118.870 105.320 119.220 106.570 ;
        RECT 122.570 105.000 122.910 105.830 ;
        RECT 124.390 105.320 124.740 106.570 ;
        RECT 128.090 105.000 128.430 105.830 ;
        RECT 129.910 105.320 130.260 106.570 ;
        RECT 133.610 105.000 133.950 105.830 ;
        RECT 135.430 105.320 135.780 106.570 ;
        RECT 138.005 105.915 139.215 107.005 ;
        RECT 138.005 105.375 138.525 105.915 ;
        RECT 138.695 105.205 139.215 105.745 ;
        RECT 115.465 104.455 120.810 105.000 ;
        RECT 120.985 104.455 126.330 105.000 ;
        RECT 126.505 104.455 131.850 105.000 ;
        RECT 132.025 104.455 137.370 105.000 ;
        RECT 138.005 104.455 139.215 105.205 ;
        RECT 50.520 104.285 139.300 104.455 ;
        RECT 50.605 103.535 51.815 104.285 ;
        RECT 52.075 103.735 52.245 104.115 ;
        RECT 52.425 103.905 52.755 104.285 ;
        RECT 52.075 103.565 52.740 103.735 ;
        RECT 52.935 103.610 53.195 104.115 ;
        RECT 53.365 103.740 58.710 104.285 ;
        RECT 50.605 102.995 51.125 103.535 ;
        RECT 51.295 102.825 51.815 103.365 ;
        RECT 52.005 103.015 52.345 103.385 ;
        RECT 52.570 103.310 52.740 103.565 ;
        RECT 52.570 102.980 52.845 103.310 ;
        RECT 52.570 102.835 52.740 102.980 ;
        RECT 50.605 101.735 51.815 102.825 ;
        RECT 52.065 102.665 52.740 102.835 ;
        RECT 53.015 102.810 53.195 103.610 ;
        RECT 54.950 102.910 55.290 103.740 ;
        RECT 59.805 103.655 60.145 104.115 ;
        RECT 60.315 103.825 60.485 104.285 ;
        RECT 60.655 103.905 61.825 104.115 ;
        RECT 60.655 103.655 60.905 103.905 ;
        RECT 61.495 103.885 61.825 103.905 ;
        RECT 62.105 103.755 62.365 104.090 ;
        RECT 62.535 103.775 62.870 104.285 ;
        RECT 63.040 103.775 63.750 104.115 ;
        RECT 59.805 103.485 60.905 103.655 ;
        RECT 61.075 103.465 61.935 103.715 ;
        RECT 52.065 101.905 52.245 102.665 ;
        RECT 52.425 101.735 52.755 102.495 ;
        RECT 52.925 101.905 53.195 102.810 ;
        RECT 56.770 102.170 57.120 103.420 ;
        RECT 59.805 103.045 60.565 103.295 ;
        RECT 60.735 103.045 61.485 103.295 ;
        RECT 61.655 102.875 61.935 103.465 ;
        RECT 53.365 101.735 58.710 102.170 ;
        RECT 59.805 101.735 60.065 102.875 ;
        RECT 60.235 102.705 61.935 102.875 ;
        RECT 60.235 101.905 60.565 102.705 ;
        RECT 60.735 101.735 60.905 102.535 ;
        RECT 61.075 101.905 61.405 102.705 ;
        RECT 61.575 101.735 61.830 102.535 ;
        RECT 62.105 102.525 62.340 103.755 ;
        RECT 62.510 102.695 62.800 103.605 ;
        RECT 62.970 103.095 63.300 103.605 ;
        RECT 63.470 103.345 63.750 103.775 ;
        RECT 63.920 103.715 64.190 104.115 ;
        RECT 64.360 103.885 64.690 104.285 ;
        RECT 64.860 103.905 66.070 104.095 ;
        RECT 64.860 103.715 65.145 103.905 ;
        RECT 66.245 103.740 71.590 104.285 ;
        RECT 63.920 103.515 65.145 103.715 ;
        RECT 65.315 103.515 66.075 103.735 ;
        RECT 63.470 103.095 64.985 103.345 ;
        RECT 65.265 103.095 65.675 103.345 ;
        RECT 63.470 102.925 63.755 103.095 ;
        RECT 65.845 102.925 66.075 103.515 ;
        RECT 63.140 102.605 63.755 102.925 ;
        RECT 63.925 102.745 66.075 102.925 ;
        RECT 67.830 102.910 68.170 103.740 ;
        RECT 71.765 103.515 75.275 104.285 ;
        RECT 76.365 103.560 76.655 104.285 ;
        RECT 76.825 103.740 82.170 104.285 ;
        RECT 82.345 103.740 87.690 104.285 ;
        RECT 87.865 103.740 93.210 104.285 ;
        RECT 93.385 103.740 98.730 104.285 ;
        RECT 63.925 102.605 65.645 102.745 ;
        RECT 62.105 101.905 62.365 102.525 ;
        RECT 62.535 101.735 62.970 102.525 ;
        RECT 63.140 101.905 63.430 102.605 ;
        RECT 63.620 102.265 65.145 102.435 ;
        RECT 63.620 101.905 63.830 102.265 ;
        RECT 64.000 101.735 64.330 102.095 ;
        RECT 64.500 102.075 65.145 102.265 ;
        RECT 65.315 102.245 65.645 102.605 ;
        RECT 65.815 102.075 66.075 102.575 ;
        RECT 69.650 102.170 70.000 103.420 ;
        RECT 71.765 102.995 73.415 103.515 ;
        RECT 73.585 102.825 75.275 103.345 ;
        RECT 78.410 102.910 78.750 103.740 ;
        RECT 64.500 101.905 66.075 102.075 ;
        RECT 66.245 101.735 71.590 102.170 ;
        RECT 71.765 101.735 75.275 102.825 ;
        RECT 76.365 101.735 76.655 102.900 ;
        RECT 80.230 102.170 80.580 103.420 ;
        RECT 83.930 102.910 84.270 103.740 ;
        RECT 85.750 102.170 86.100 103.420 ;
        RECT 89.450 102.910 89.790 103.740 ;
        RECT 91.270 102.170 91.620 103.420 ;
        RECT 94.970 102.910 95.310 103.740 ;
        RECT 98.905 103.515 101.495 104.285 ;
        RECT 102.125 103.560 102.415 104.285 ;
        RECT 102.585 103.740 107.930 104.285 ;
        RECT 108.105 103.740 113.450 104.285 ;
        RECT 113.625 103.740 118.970 104.285 ;
        RECT 119.145 103.740 124.490 104.285 ;
        RECT 96.790 102.170 97.140 103.420 ;
        RECT 98.905 102.995 100.115 103.515 ;
        RECT 100.285 102.825 101.495 103.345 ;
        RECT 104.170 102.910 104.510 103.740 ;
        RECT 76.825 101.735 82.170 102.170 ;
        RECT 82.345 101.735 87.690 102.170 ;
        RECT 87.865 101.735 93.210 102.170 ;
        RECT 93.385 101.735 98.730 102.170 ;
        RECT 98.905 101.735 101.495 102.825 ;
        RECT 102.125 101.735 102.415 102.900 ;
        RECT 105.990 102.170 106.340 103.420 ;
        RECT 109.690 102.910 110.030 103.740 ;
        RECT 111.510 102.170 111.860 103.420 ;
        RECT 115.210 102.910 115.550 103.740 ;
        RECT 117.030 102.170 117.380 103.420 ;
        RECT 120.730 102.910 121.070 103.740 ;
        RECT 124.665 103.515 127.255 104.285 ;
        RECT 127.885 103.560 128.175 104.285 ;
        RECT 128.345 103.740 133.690 104.285 ;
        RECT 122.550 102.170 122.900 103.420 ;
        RECT 124.665 102.995 125.875 103.515 ;
        RECT 126.045 102.825 127.255 103.345 ;
        RECT 129.930 102.910 130.270 103.740 ;
        RECT 133.865 103.515 137.375 104.285 ;
        RECT 138.005 103.535 139.215 104.285 ;
        RECT 102.585 101.735 107.930 102.170 ;
        RECT 108.105 101.735 113.450 102.170 ;
        RECT 113.625 101.735 118.970 102.170 ;
        RECT 119.145 101.735 124.490 102.170 ;
        RECT 124.665 101.735 127.255 102.825 ;
        RECT 127.885 101.735 128.175 102.900 ;
        RECT 131.750 102.170 132.100 103.420 ;
        RECT 133.865 102.995 135.515 103.515 ;
        RECT 135.685 102.825 137.375 103.345 ;
        RECT 128.345 101.735 133.690 102.170 ;
        RECT 133.865 101.735 137.375 102.825 ;
        RECT 138.005 102.825 138.525 103.365 ;
        RECT 138.695 102.995 139.215 103.535 ;
        RECT 138.005 101.735 139.215 102.825 ;
        RECT 50.520 101.565 139.300 101.735 ;
        RECT 50.605 100.475 51.815 101.565 ;
        RECT 50.605 99.765 51.125 100.305 ;
        RECT 51.295 99.935 51.815 100.475 ;
        RECT 52.065 100.635 52.245 101.395 ;
        RECT 52.425 100.805 52.755 101.565 ;
        RECT 52.065 100.465 52.740 100.635 ;
        RECT 52.925 100.490 53.195 101.395 ;
        RECT 53.365 101.130 58.710 101.565 ;
        RECT 52.570 100.320 52.740 100.465 ;
        RECT 52.005 99.915 52.345 100.285 ;
        RECT 52.570 99.990 52.845 100.320 ;
        RECT 50.605 99.015 51.815 99.765 ;
        RECT 52.570 99.735 52.740 99.990 ;
        RECT 52.075 99.565 52.740 99.735 ;
        RECT 53.015 99.690 53.195 100.490 ;
        RECT 52.075 99.185 52.245 99.565 ;
        RECT 52.425 99.015 52.755 99.395 ;
        RECT 52.935 99.185 53.195 99.690 ;
        RECT 54.950 99.560 55.290 100.390 ;
        RECT 56.770 99.880 57.120 101.130 ;
        RECT 58.885 100.475 62.395 101.565 ;
        RECT 58.885 99.785 60.535 100.305 ;
        RECT 60.705 99.955 62.395 100.475 ;
        RECT 63.485 100.400 63.775 101.565 ;
        RECT 63.945 101.130 69.290 101.565 ;
        RECT 69.465 101.130 74.810 101.565 ;
        RECT 74.985 101.130 80.330 101.565 ;
        RECT 80.505 101.130 85.850 101.565 ;
        RECT 53.365 99.015 58.710 99.560 ;
        RECT 58.885 99.015 62.395 99.785 ;
        RECT 63.485 99.015 63.775 99.740 ;
        RECT 65.530 99.560 65.870 100.390 ;
        RECT 67.350 99.880 67.700 101.130 ;
        RECT 71.050 99.560 71.390 100.390 ;
        RECT 72.870 99.880 73.220 101.130 ;
        RECT 76.570 99.560 76.910 100.390 ;
        RECT 78.390 99.880 78.740 101.130 ;
        RECT 82.090 99.560 82.430 100.390 ;
        RECT 83.910 99.880 84.260 101.130 ;
        RECT 86.025 100.475 88.615 101.565 ;
        RECT 86.025 99.785 87.235 100.305 ;
        RECT 87.405 99.955 88.615 100.475 ;
        RECT 89.245 100.400 89.535 101.565 ;
        RECT 89.705 101.130 95.050 101.565 ;
        RECT 95.225 101.130 100.570 101.565 ;
        RECT 100.745 101.130 106.090 101.565 ;
        RECT 106.265 101.130 111.610 101.565 ;
        RECT 63.945 99.015 69.290 99.560 ;
        RECT 69.465 99.015 74.810 99.560 ;
        RECT 74.985 99.015 80.330 99.560 ;
        RECT 80.505 99.015 85.850 99.560 ;
        RECT 86.025 99.015 88.615 99.785 ;
        RECT 89.245 99.015 89.535 99.740 ;
        RECT 91.290 99.560 91.630 100.390 ;
        RECT 93.110 99.880 93.460 101.130 ;
        RECT 96.810 99.560 97.150 100.390 ;
        RECT 98.630 99.880 98.980 101.130 ;
        RECT 102.330 99.560 102.670 100.390 ;
        RECT 104.150 99.880 104.500 101.130 ;
        RECT 107.850 99.560 108.190 100.390 ;
        RECT 109.670 99.880 110.020 101.130 ;
        RECT 111.785 100.475 114.375 101.565 ;
        RECT 111.785 99.785 112.995 100.305 ;
        RECT 113.165 99.955 114.375 100.475 ;
        RECT 115.005 100.400 115.295 101.565 ;
        RECT 115.465 101.130 120.810 101.565 ;
        RECT 120.985 101.130 126.330 101.565 ;
        RECT 126.505 101.130 131.850 101.565 ;
        RECT 132.025 101.130 137.370 101.565 ;
        RECT 89.705 99.015 95.050 99.560 ;
        RECT 95.225 99.015 100.570 99.560 ;
        RECT 100.745 99.015 106.090 99.560 ;
        RECT 106.265 99.015 111.610 99.560 ;
        RECT 111.785 99.015 114.375 99.785 ;
        RECT 115.005 99.015 115.295 99.740 ;
        RECT 117.050 99.560 117.390 100.390 ;
        RECT 118.870 99.880 119.220 101.130 ;
        RECT 122.570 99.560 122.910 100.390 ;
        RECT 124.390 99.880 124.740 101.130 ;
        RECT 128.090 99.560 128.430 100.390 ;
        RECT 129.910 99.880 130.260 101.130 ;
        RECT 133.610 99.560 133.950 100.390 ;
        RECT 135.430 99.880 135.780 101.130 ;
        RECT 138.005 100.475 139.215 101.565 ;
        RECT 138.005 99.935 138.525 100.475 ;
        RECT 138.695 99.765 139.215 100.305 ;
        RECT 115.465 99.015 120.810 99.560 ;
        RECT 120.985 99.015 126.330 99.560 ;
        RECT 126.505 99.015 131.850 99.560 ;
        RECT 132.025 99.015 137.370 99.560 ;
        RECT 138.005 99.015 139.215 99.765 ;
        RECT 50.520 98.845 139.300 99.015 ;
        RECT 50.605 98.095 51.815 98.845 ;
        RECT 51.985 98.300 57.330 98.845 ;
        RECT 50.605 97.555 51.125 98.095 ;
        RECT 51.295 97.385 51.815 97.925 ;
        RECT 53.570 97.470 53.910 98.300 ;
        RECT 57.505 98.075 60.095 98.845 ;
        RECT 60.815 98.295 60.985 98.675 ;
        RECT 61.165 98.465 61.495 98.845 ;
        RECT 60.815 98.125 61.480 98.295 ;
        RECT 61.675 98.170 61.935 98.675 ;
        RECT 62.105 98.300 67.450 98.845 ;
        RECT 67.625 98.300 72.970 98.845 ;
        RECT 50.605 96.295 51.815 97.385 ;
        RECT 55.390 96.730 55.740 97.980 ;
        RECT 57.505 97.555 58.715 98.075 ;
        RECT 58.885 97.385 60.095 97.905 ;
        RECT 60.745 97.575 61.075 97.945 ;
        RECT 61.310 97.870 61.480 98.125 ;
        RECT 61.310 97.540 61.595 97.870 ;
        RECT 61.310 97.395 61.480 97.540 ;
        RECT 51.985 96.295 57.330 96.730 ;
        RECT 57.505 96.295 60.095 97.385 ;
        RECT 60.815 97.225 61.480 97.395 ;
        RECT 61.765 97.370 61.935 98.170 ;
        RECT 63.690 97.470 64.030 98.300 ;
        RECT 60.815 96.465 60.985 97.225 ;
        RECT 61.165 96.295 61.495 97.055 ;
        RECT 61.665 96.465 61.935 97.370 ;
        RECT 65.510 96.730 65.860 97.980 ;
        RECT 69.210 97.470 69.550 98.300 ;
        RECT 73.145 98.075 75.735 98.845 ;
        RECT 76.365 98.120 76.655 98.845 ;
        RECT 76.825 98.300 82.170 98.845 ;
        RECT 82.345 98.300 87.690 98.845 ;
        RECT 87.865 98.300 93.210 98.845 ;
        RECT 93.385 98.300 98.730 98.845 ;
        RECT 71.030 96.730 71.380 97.980 ;
        RECT 73.145 97.555 74.355 98.075 ;
        RECT 74.525 97.385 75.735 97.905 ;
        RECT 78.410 97.470 78.750 98.300 ;
        RECT 62.105 96.295 67.450 96.730 ;
        RECT 67.625 96.295 72.970 96.730 ;
        RECT 73.145 96.295 75.735 97.385 ;
        RECT 76.365 96.295 76.655 97.460 ;
        RECT 80.230 96.730 80.580 97.980 ;
        RECT 83.930 97.470 84.270 98.300 ;
        RECT 85.750 96.730 86.100 97.980 ;
        RECT 89.450 97.470 89.790 98.300 ;
        RECT 91.270 96.730 91.620 97.980 ;
        RECT 94.970 97.470 95.310 98.300 ;
        RECT 98.905 98.075 101.495 98.845 ;
        RECT 102.125 98.120 102.415 98.845 ;
        RECT 102.585 98.300 107.930 98.845 ;
        RECT 108.105 98.300 113.450 98.845 ;
        RECT 113.625 98.300 118.970 98.845 ;
        RECT 119.145 98.300 124.490 98.845 ;
        RECT 96.790 96.730 97.140 97.980 ;
        RECT 98.905 97.555 100.115 98.075 ;
        RECT 100.285 97.385 101.495 97.905 ;
        RECT 104.170 97.470 104.510 98.300 ;
        RECT 76.825 96.295 82.170 96.730 ;
        RECT 82.345 96.295 87.690 96.730 ;
        RECT 87.865 96.295 93.210 96.730 ;
        RECT 93.385 96.295 98.730 96.730 ;
        RECT 98.905 96.295 101.495 97.385 ;
        RECT 102.125 96.295 102.415 97.460 ;
        RECT 105.990 96.730 106.340 97.980 ;
        RECT 109.690 97.470 110.030 98.300 ;
        RECT 111.510 96.730 111.860 97.980 ;
        RECT 115.210 97.470 115.550 98.300 ;
        RECT 117.030 96.730 117.380 97.980 ;
        RECT 120.730 97.470 121.070 98.300 ;
        RECT 124.665 98.075 127.255 98.845 ;
        RECT 127.885 98.120 128.175 98.845 ;
        RECT 128.345 98.300 133.690 98.845 ;
        RECT 122.550 96.730 122.900 97.980 ;
        RECT 124.665 97.555 125.875 98.075 ;
        RECT 126.045 97.385 127.255 97.905 ;
        RECT 129.930 97.470 130.270 98.300 ;
        RECT 133.865 98.075 137.375 98.845 ;
        RECT 138.005 98.095 139.215 98.845 ;
        RECT 102.585 96.295 107.930 96.730 ;
        RECT 108.105 96.295 113.450 96.730 ;
        RECT 113.625 96.295 118.970 96.730 ;
        RECT 119.145 96.295 124.490 96.730 ;
        RECT 124.665 96.295 127.255 97.385 ;
        RECT 127.885 96.295 128.175 97.460 ;
        RECT 131.750 96.730 132.100 97.980 ;
        RECT 133.865 97.555 135.515 98.075 ;
        RECT 135.685 97.385 137.375 97.905 ;
        RECT 128.345 96.295 133.690 96.730 ;
        RECT 133.865 96.295 137.375 97.385 ;
        RECT 138.005 97.385 138.525 97.925 ;
        RECT 138.695 97.555 139.215 98.095 ;
        RECT 138.005 96.295 139.215 97.385 ;
        RECT 50.520 96.125 139.300 96.295 ;
        RECT 50.605 95.035 51.815 96.125 ;
        RECT 51.985 95.690 57.330 96.125 ;
        RECT 50.605 94.325 51.125 94.865 ;
        RECT 51.295 94.495 51.815 95.035 ;
        RECT 50.605 93.575 51.815 94.325 ;
        RECT 53.570 94.120 53.910 94.950 ;
        RECT 55.390 94.440 55.740 95.690 ;
        RECT 57.505 95.035 61.015 96.125 ;
        RECT 57.505 94.345 59.155 94.865 ;
        RECT 59.325 94.515 61.015 95.035 ;
        RECT 61.645 94.985 61.905 96.125 ;
        RECT 62.075 94.975 62.405 95.955 ;
        RECT 62.575 94.985 62.855 96.125 ;
        RECT 61.665 94.565 62.000 94.815 ;
        RECT 62.170 94.375 62.340 94.975 ;
        RECT 63.485 94.960 63.775 96.125 ;
        RECT 63.945 95.690 69.290 96.125 ;
        RECT 69.465 95.690 74.810 96.125 ;
        RECT 74.985 95.690 80.330 96.125 ;
        RECT 80.505 95.690 85.850 96.125 ;
        RECT 62.510 94.545 62.845 94.815 ;
        RECT 51.985 93.575 57.330 94.120 ;
        RECT 57.505 93.575 61.015 94.345 ;
        RECT 61.645 93.745 62.340 94.375 ;
        RECT 62.545 93.575 62.855 94.375 ;
        RECT 63.485 93.575 63.775 94.300 ;
        RECT 65.530 94.120 65.870 94.950 ;
        RECT 67.350 94.440 67.700 95.690 ;
        RECT 71.050 94.120 71.390 94.950 ;
        RECT 72.870 94.440 73.220 95.690 ;
        RECT 76.570 94.120 76.910 94.950 ;
        RECT 78.390 94.440 78.740 95.690 ;
        RECT 82.090 94.120 82.430 94.950 ;
        RECT 83.910 94.440 84.260 95.690 ;
        RECT 86.025 95.035 88.615 96.125 ;
        RECT 86.025 94.345 87.235 94.865 ;
        RECT 87.405 94.515 88.615 95.035 ;
        RECT 89.245 94.960 89.535 96.125 ;
        RECT 89.705 95.690 95.050 96.125 ;
        RECT 95.225 95.690 100.570 96.125 ;
        RECT 100.745 95.690 106.090 96.125 ;
        RECT 106.265 95.690 111.610 96.125 ;
        RECT 63.945 93.575 69.290 94.120 ;
        RECT 69.465 93.575 74.810 94.120 ;
        RECT 74.985 93.575 80.330 94.120 ;
        RECT 80.505 93.575 85.850 94.120 ;
        RECT 86.025 93.575 88.615 94.345 ;
        RECT 89.245 93.575 89.535 94.300 ;
        RECT 91.290 94.120 91.630 94.950 ;
        RECT 93.110 94.440 93.460 95.690 ;
        RECT 96.810 94.120 97.150 94.950 ;
        RECT 98.630 94.440 98.980 95.690 ;
        RECT 102.330 94.120 102.670 94.950 ;
        RECT 104.150 94.440 104.500 95.690 ;
        RECT 107.850 94.120 108.190 94.950 ;
        RECT 109.670 94.440 110.020 95.690 ;
        RECT 111.785 95.035 114.375 96.125 ;
        RECT 111.785 94.345 112.995 94.865 ;
        RECT 113.165 94.515 114.375 95.035 ;
        RECT 115.005 94.960 115.295 96.125 ;
        RECT 115.465 95.690 120.810 96.125 ;
        RECT 120.985 95.690 126.330 96.125 ;
        RECT 126.505 95.690 131.850 96.125 ;
        RECT 132.025 95.690 137.370 96.125 ;
        RECT 89.705 93.575 95.050 94.120 ;
        RECT 95.225 93.575 100.570 94.120 ;
        RECT 100.745 93.575 106.090 94.120 ;
        RECT 106.265 93.575 111.610 94.120 ;
        RECT 111.785 93.575 114.375 94.345 ;
        RECT 115.005 93.575 115.295 94.300 ;
        RECT 117.050 94.120 117.390 94.950 ;
        RECT 118.870 94.440 119.220 95.690 ;
        RECT 122.570 94.120 122.910 94.950 ;
        RECT 124.390 94.440 124.740 95.690 ;
        RECT 128.090 94.120 128.430 94.950 ;
        RECT 129.910 94.440 130.260 95.690 ;
        RECT 133.610 94.120 133.950 94.950 ;
        RECT 135.430 94.440 135.780 95.690 ;
        RECT 138.005 95.035 139.215 96.125 ;
        RECT 138.005 94.495 138.525 95.035 ;
        RECT 138.695 94.325 139.215 94.865 ;
        RECT 115.465 93.575 120.810 94.120 ;
        RECT 120.985 93.575 126.330 94.120 ;
        RECT 126.505 93.575 131.850 94.120 ;
        RECT 132.025 93.575 137.370 94.120 ;
        RECT 138.005 93.575 139.215 94.325 ;
        RECT 50.520 93.405 139.300 93.575 ;
        RECT 50.605 92.655 51.815 93.405 ;
        RECT 50.605 92.115 51.125 92.655 ;
        RECT 51.985 92.635 55.495 93.405 ;
        RECT 51.295 91.945 51.815 92.485 ;
        RECT 51.985 92.115 53.635 92.635 ;
        RECT 56.860 92.595 57.105 93.200 ;
        RECT 57.325 92.870 57.835 93.405 ;
        RECT 53.805 91.945 55.495 92.465 ;
        RECT 50.605 90.855 51.815 91.945 ;
        RECT 51.985 90.855 55.495 91.945 ;
        RECT 56.585 92.425 57.815 92.595 ;
        RECT 56.585 91.615 56.925 92.425 ;
        RECT 57.095 91.860 57.845 92.050 ;
        RECT 56.585 91.205 57.100 91.615 ;
        RECT 57.335 90.855 57.505 91.615 ;
        RECT 57.675 91.195 57.845 91.860 ;
        RECT 58.015 91.875 58.205 93.235 ;
        RECT 58.375 93.065 58.650 93.235 ;
        RECT 58.375 92.895 58.655 93.065 ;
        RECT 58.375 92.075 58.650 92.895 ;
        RECT 58.840 92.870 59.370 93.235 ;
        RECT 59.795 93.005 60.125 93.405 ;
        RECT 59.195 92.835 59.370 92.870 ;
        RECT 58.855 91.875 59.025 92.675 ;
        RECT 58.015 91.705 59.025 91.875 ;
        RECT 59.195 92.665 60.125 92.835 ;
        RECT 60.295 92.665 60.550 93.235 ;
        RECT 59.195 91.535 59.365 92.665 ;
        RECT 59.955 92.495 60.125 92.665 ;
        RECT 58.240 91.365 59.365 91.535 ;
        RECT 59.535 92.165 59.730 92.495 ;
        RECT 59.955 92.165 60.210 92.495 ;
        RECT 59.535 91.195 59.705 92.165 ;
        RECT 60.380 91.995 60.550 92.665 ;
        RECT 57.675 91.025 59.705 91.195 ;
        RECT 59.875 90.855 60.045 91.995 ;
        RECT 60.215 91.025 60.550 91.995 ;
        RECT 60.730 92.665 60.985 93.235 ;
        RECT 61.155 93.005 61.485 93.405 ;
        RECT 61.910 92.870 62.440 93.235 ;
        RECT 61.910 92.835 62.085 92.870 ;
        RECT 61.155 92.665 62.085 92.835 ;
        RECT 60.730 91.995 60.900 92.665 ;
        RECT 61.155 92.495 61.325 92.665 ;
        RECT 61.070 92.165 61.325 92.495 ;
        RECT 61.550 92.165 61.745 92.495 ;
        RECT 60.730 91.025 61.065 91.995 ;
        RECT 61.235 90.855 61.405 91.995 ;
        RECT 61.575 91.195 61.745 92.165 ;
        RECT 61.915 91.535 62.085 92.665 ;
        RECT 62.255 91.875 62.425 92.675 ;
        RECT 62.630 92.385 62.905 93.235 ;
        RECT 62.625 92.215 62.905 92.385 ;
        RECT 62.630 92.075 62.905 92.215 ;
        RECT 63.075 91.875 63.265 93.235 ;
        RECT 63.445 92.870 63.955 93.405 ;
        RECT 64.175 92.595 64.420 93.200 ;
        RECT 63.465 92.425 64.695 92.595 ;
        RECT 64.905 92.585 65.135 93.405 ;
        RECT 65.305 92.605 65.635 93.235 ;
        RECT 62.255 91.705 63.265 91.875 ;
        RECT 63.435 91.860 64.185 92.050 ;
        RECT 61.915 91.365 63.040 91.535 ;
        RECT 63.435 91.195 63.605 91.860 ;
        RECT 64.355 91.615 64.695 92.425 ;
        RECT 64.885 92.165 65.215 92.415 ;
        RECT 65.385 92.005 65.635 92.605 ;
        RECT 65.805 92.585 66.015 93.405 ;
        RECT 66.285 92.585 66.515 93.405 ;
        RECT 66.685 92.605 67.015 93.235 ;
        RECT 66.265 92.165 66.595 92.415 ;
        RECT 66.765 92.005 67.015 92.605 ;
        RECT 67.185 92.585 67.395 93.405 ;
        RECT 67.625 92.860 72.970 93.405 ;
        RECT 69.210 92.030 69.550 92.860 ;
        RECT 73.145 92.635 75.735 93.405 ;
        RECT 76.365 92.680 76.655 93.405 ;
        RECT 76.825 92.860 82.170 93.405 ;
        RECT 82.345 92.860 87.690 93.405 ;
        RECT 87.865 92.860 93.210 93.405 ;
        RECT 93.385 92.860 98.730 93.405 ;
        RECT 61.575 91.025 63.605 91.195 ;
        RECT 63.775 90.855 63.945 91.615 ;
        RECT 64.180 91.205 64.695 91.615 ;
        RECT 64.905 90.855 65.135 91.995 ;
        RECT 65.305 91.025 65.635 92.005 ;
        RECT 65.805 90.855 66.015 91.995 ;
        RECT 66.285 90.855 66.515 91.995 ;
        RECT 66.685 91.025 67.015 92.005 ;
        RECT 67.185 90.855 67.395 91.995 ;
        RECT 71.030 91.290 71.380 92.540 ;
        RECT 73.145 92.115 74.355 92.635 ;
        RECT 74.525 91.945 75.735 92.465 ;
        RECT 78.410 92.030 78.750 92.860 ;
        RECT 67.625 90.855 72.970 91.290 ;
        RECT 73.145 90.855 75.735 91.945 ;
        RECT 76.365 90.855 76.655 92.020 ;
        RECT 80.230 91.290 80.580 92.540 ;
        RECT 83.930 92.030 84.270 92.860 ;
        RECT 85.750 91.290 86.100 92.540 ;
        RECT 89.450 92.030 89.790 92.860 ;
        RECT 91.270 91.290 91.620 92.540 ;
        RECT 94.970 92.030 95.310 92.860 ;
        RECT 98.905 92.635 101.495 93.405 ;
        RECT 102.125 92.680 102.415 93.405 ;
        RECT 102.585 92.860 107.930 93.405 ;
        RECT 108.105 92.860 113.450 93.405 ;
        RECT 113.625 92.860 118.970 93.405 ;
        RECT 119.145 92.860 124.490 93.405 ;
        RECT 96.790 91.290 97.140 92.540 ;
        RECT 98.905 92.115 100.115 92.635 ;
        RECT 100.285 91.945 101.495 92.465 ;
        RECT 104.170 92.030 104.510 92.860 ;
        RECT 76.825 90.855 82.170 91.290 ;
        RECT 82.345 90.855 87.690 91.290 ;
        RECT 87.865 90.855 93.210 91.290 ;
        RECT 93.385 90.855 98.730 91.290 ;
        RECT 98.905 90.855 101.495 91.945 ;
        RECT 102.125 90.855 102.415 92.020 ;
        RECT 105.990 91.290 106.340 92.540 ;
        RECT 109.690 92.030 110.030 92.860 ;
        RECT 111.510 91.290 111.860 92.540 ;
        RECT 115.210 92.030 115.550 92.860 ;
        RECT 117.030 91.290 117.380 92.540 ;
        RECT 120.730 92.030 121.070 92.860 ;
        RECT 124.665 92.635 127.255 93.405 ;
        RECT 127.885 92.680 128.175 93.405 ;
        RECT 128.345 92.860 133.690 93.405 ;
        RECT 122.550 91.290 122.900 92.540 ;
        RECT 124.665 92.115 125.875 92.635 ;
        RECT 126.045 91.945 127.255 92.465 ;
        RECT 129.930 92.030 130.270 92.860 ;
        RECT 133.865 92.635 137.375 93.405 ;
        RECT 138.005 92.655 139.215 93.405 ;
        RECT 102.585 90.855 107.930 91.290 ;
        RECT 108.105 90.855 113.450 91.290 ;
        RECT 113.625 90.855 118.970 91.290 ;
        RECT 119.145 90.855 124.490 91.290 ;
        RECT 124.665 90.855 127.255 91.945 ;
        RECT 127.885 90.855 128.175 92.020 ;
        RECT 131.750 91.290 132.100 92.540 ;
        RECT 133.865 92.115 135.515 92.635 ;
        RECT 135.685 91.945 137.375 92.465 ;
        RECT 128.345 90.855 133.690 91.290 ;
        RECT 133.865 90.855 137.375 91.945 ;
        RECT 138.005 91.945 138.525 92.485 ;
        RECT 138.695 92.115 139.215 92.655 ;
        RECT 138.005 90.855 139.215 91.945 ;
        RECT 50.520 90.685 139.300 90.855 ;
        RECT 50.605 89.595 51.815 90.685 ;
        RECT 51.985 90.250 57.330 90.685 ;
        RECT 50.605 88.885 51.125 89.425 ;
        RECT 51.295 89.055 51.815 89.595 ;
        RECT 50.605 88.135 51.815 88.885 ;
        RECT 53.570 88.680 53.910 89.510 ;
        RECT 55.390 89.000 55.740 90.250 ;
        RECT 57.505 89.595 60.095 90.685 ;
        RECT 57.505 88.905 58.715 89.425 ;
        RECT 58.885 89.075 60.095 89.595 ;
        RECT 60.345 89.755 60.525 90.515 ;
        RECT 60.705 89.925 61.035 90.685 ;
        RECT 60.345 89.585 61.020 89.755 ;
        RECT 61.205 89.610 61.475 90.515 ;
        RECT 60.850 89.440 61.020 89.585 ;
        RECT 60.285 89.035 60.625 89.405 ;
        RECT 60.850 89.110 61.125 89.440 ;
        RECT 51.985 88.135 57.330 88.680 ;
        RECT 57.505 88.135 60.095 88.905 ;
        RECT 60.850 88.855 61.020 89.110 ;
        RECT 60.355 88.685 61.020 88.855 ;
        RECT 61.295 88.810 61.475 89.610 ;
        RECT 61.685 89.545 61.915 90.685 ;
        RECT 62.085 89.535 62.415 90.515 ;
        RECT 62.585 89.545 62.795 90.685 ;
        RECT 61.665 89.125 61.995 89.375 ;
        RECT 60.355 88.305 60.525 88.685 ;
        RECT 60.705 88.135 61.035 88.515 ;
        RECT 61.215 88.305 61.475 88.810 ;
        RECT 61.685 88.135 61.915 88.955 ;
        RECT 62.165 88.935 62.415 89.535 ;
        RECT 63.485 89.520 63.775 90.685 ;
        RECT 63.945 90.250 69.290 90.685 ;
        RECT 69.465 90.250 74.810 90.685 ;
        RECT 74.985 90.250 80.330 90.685 ;
        RECT 80.505 90.250 85.850 90.685 ;
        RECT 62.085 88.305 62.415 88.935 ;
        RECT 62.585 88.135 62.795 88.955 ;
        RECT 63.485 88.135 63.775 88.860 ;
        RECT 65.530 88.680 65.870 89.510 ;
        RECT 67.350 89.000 67.700 90.250 ;
        RECT 71.050 88.680 71.390 89.510 ;
        RECT 72.870 89.000 73.220 90.250 ;
        RECT 76.570 88.680 76.910 89.510 ;
        RECT 78.390 89.000 78.740 90.250 ;
        RECT 82.090 88.680 82.430 89.510 ;
        RECT 83.910 89.000 84.260 90.250 ;
        RECT 86.025 89.595 88.615 90.685 ;
        RECT 86.025 88.905 87.235 89.425 ;
        RECT 87.405 89.075 88.615 89.595 ;
        RECT 89.245 89.520 89.535 90.685 ;
        RECT 89.705 90.250 95.050 90.685 ;
        RECT 95.225 90.250 100.570 90.685 ;
        RECT 100.745 90.250 106.090 90.685 ;
        RECT 106.265 90.250 111.610 90.685 ;
        RECT 63.945 88.135 69.290 88.680 ;
        RECT 69.465 88.135 74.810 88.680 ;
        RECT 74.985 88.135 80.330 88.680 ;
        RECT 80.505 88.135 85.850 88.680 ;
        RECT 86.025 88.135 88.615 88.905 ;
        RECT 89.245 88.135 89.535 88.860 ;
        RECT 91.290 88.680 91.630 89.510 ;
        RECT 93.110 89.000 93.460 90.250 ;
        RECT 96.810 88.680 97.150 89.510 ;
        RECT 98.630 89.000 98.980 90.250 ;
        RECT 102.330 88.680 102.670 89.510 ;
        RECT 104.150 89.000 104.500 90.250 ;
        RECT 107.850 88.680 108.190 89.510 ;
        RECT 109.670 89.000 110.020 90.250 ;
        RECT 111.785 89.595 114.375 90.685 ;
        RECT 111.785 88.905 112.995 89.425 ;
        RECT 113.165 89.075 114.375 89.595 ;
        RECT 115.005 89.520 115.295 90.685 ;
        RECT 115.465 90.250 120.810 90.685 ;
        RECT 120.985 90.250 126.330 90.685 ;
        RECT 126.505 90.250 131.850 90.685 ;
        RECT 132.025 90.250 137.370 90.685 ;
        RECT 89.705 88.135 95.050 88.680 ;
        RECT 95.225 88.135 100.570 88.680 ;
        RECT 100.745 88.135 106.090 88.680 ;
        RECT 106.265 88.135 111.610 88.680 ;
        RECT 111.785 88.135 114.375 88.905 ;
        RECT 115.005 88.135 115.295 88.860 ;
        RECT 117.050 88.680 117.390 89.510 ;
        RECT 118.870 89.000 119.220 90.250 ;
        RECT 122.570 88.680 122.910 89.510 ;
        RECT 124.390 89.000 124.740 90.250 ;
        RECT 128.090 88.680 128.430 89.510 ;
        RECT 129.910 89.000 130.260 90.250 ;
        RECT 133.610 88.680 133.950 89.510 ;
        RECT 135.430 89.000 135.780 90.250 ;
        RECT 138.005 89.595 139.215 90.685 ;
        RECT 138.005 89.055 138.525 89.595 ;
        RECT 138.695 88.885 139.215 89.425 ;
        RECT 115.465 88.135 120.810 88.680 ;
        RECT 120.985 88.135 126.330 88.680 ;
        RECT 126.505 88.135 131.850 88.680 ;
        RECT 132.025 88.135 137.370 88.680 ;
        RECT 138.005 88.135 139.215 88.885 ;
        RECT 50.520 87.965 139.300 88.135 ;
        RECT 50.605 87.215 51.815 87.965 ;
        RECT 51.985 87.420 57.330 87.965 ;
        RECT 57.505 87.420 62.850 87.965 ;
        RECT 63.025 87.420 68.370 87.965 ;
        RECT 68.545 87.420 73.890 87.965 ;
        RECT 50.605 86.675 51.125 87.215 ;
        RECT 51.295 86.505 51.815 87.045 ;
        RECT 53.570 86.590 53.910 87.420 ;
        RECT 50.605 85.415 51.815 86.505 ;
        RECT 55.390 85.850 55.740 87.100 ;
        RECT 59.090 86.590 59.430 87.420 ;
        RECT 60.910 85.850 61.260 87.100 ;
        RECT 64.610 86.590 64.950 87.420 ;
        RECT 66.430 85.850 66.780 87.100 ;
        RECT 70.130 86.590 70.470 87.420 ;
        RECT 74.065 87.195 75.735 87.965 ;
        RECT 76.365 87.240 76.655 87.965 ;
        RECT 76.825 87.420 82.170 87.965 ;
        RECT 82.345 87.420 87.690 87.965 ;
        RECT 87.865 87.420 93.210 87.965 ;
        RECT 93.385 87.420 98.730 87.965 ;
        RECT 71.950 85.850 72.300 87.100 ;
        RECT 74.065 86.675 74.815 87.195 ;
        RECT 74.985 86.505 75.735 87.025 ;
        RECT 78.410 86.590 78.750 87.420 ;
        RECT 51.985 85.415 57.330 85.850 ;
        RECT 57.505 85.415 62.850 85.850 ;
        RECT 63.025 85.415 68.370 85.850 ;
        RECT 68.545 85.415 73.890 85.850 ;
        RECT 74.065 85.415 75.735 86.505 ;
        RECT 76.365 85.415 76.655 86.580 ;
        RECT 80.230 85.850 80.580 87.100 ;
        RECT 83.930 86.590 84.270 87.420 ;
        RECT 85.750 85.850 86.100 87.100 ;
        RECT 89.450 86.590 89.790 87.420 ;
        RECT 91.270 85.850 91.620 87.100 ;
        RECT 94.970 86.590 95.310 87.420 ;
        RECT 98.905 87.195 101.495 87.965 ;
        RECT 102.125 87.240 102.415 87.965 ;
        RECT 102.585 87.420 107.930 87.965 ;
        RECT 108.105 87.420 113.450 87.965 ;
        RECT 113.625 87.420 118.970 87.965 ;
        RECT 119.145 87.420 124.490 87.965 ;
        RECT 96.790 85.850 97.140 87.100 ;
        RECT 98.905 86.675 100.115 87.195 ;
        RECT 100.285 86.505 101.495 87.025 ;
        RECT 104.170 86.590 104.510 87.420 ;
        RECT 76.825 85.415 82.170 85.850 ;
        RECT 82.345 85.415 87.690 85.850 ;
        RECT 87.865 85.415 93.210 85.850 ;
        RECT 93.385 85.415 98.730 85.850 ;
        RECT 98.905 85.415 101.495 86.505 ;
        RECT 102.125 85.415 102.415 86.580 ;
        RECT 105.990 85.850 106.340 87.100 ;
        RECT 109.690 86.590 110.030 87.420 ;
        RECT 111.510 85.850 111.860 87.100 ;
        RECT 115.210 86.590 115.550 87.420 ;
        RECT 117.030 85.850 117.380 87.100 ;
        RECT 120.730 86.590 121.070 87.420 ;
        RECT 124.665 87.195 127.255 87.965 ;
        RECT 127.885 87.240 128.175 87.965 ;
        RECT 128.345 87.420 133.690 87.965 ;
        RECT 122.550 85.850 122.900 87.100 ;
        RECT 124.665 86.675 125.875 87.195 ;
        RECT 126.045 86.505 127.255 87.025 ;
        RECT 129.930 86.590 130.270 87.420 ;
        RECT 133.865 87.195 137.375 87.965 ;
        RECT 138.005 87.215 139.215 87.965 ;
        RECT 102.585 85.415 107.930 85.850 ;
        RECT 108.105 85.415 113.450 85.850 ;
        RECT 113.625 85.415 118.970 85.850 ;
        RECT 119.145 85.415 124.490 85.850 ;
        RECT 124.665 85.415 127.255 86.505 ;
        RECT 127.885 85.415 128.175 86.580 ;
        RECT 131.750 85.850 132.100 87.100 ;
        RECT 133.865 86.675 135.515 87.195 ;
        RECT 135.685 86.505 137.375 87.025 ;
        RECT 128.345 85.415 133.690 85.850 ;
        RECT 133.865 85.415 137.375 86.505 ;
        RECT 138.005 86.505 138.525 87.045 ;
        RECT 138.695 86.675 139.215 87.215 ;
        RECT 138.005 85.415 139.215 86.505 ;
        RECT 50.520 85.245 139.300 85.415 ;
        RECT 50.605 84.155 51.815 85.245 ;
        RECT 51.985 84.810 57.330 85.245 ;
        RECT 57.505 84.810 62.850 85.245 ;
        RECT 50.605 83.445 51.125 83.985 ;
        RECT 51.295 83.615 51.815 84.155 ;
        RECT 50.605 82.695 51.815 83.445 ;
        RECT 53.570 83.240 53.910 84.070 ;
        RECT 55.390 83.560 55.740 84.810 ;
        RECT 59.090 83.240 59.430 84.070 ;
        RECT 60.910 83.560 61.260 84.810 ;
        RECT 63.485 84.080 63.775 85.245 ;
        RECT 63.945 84.810 69.290 85.245 ;
        RECT 69.465 84.810 74.810 85.245 ;
        RECT 74.985 84.810 80.330 85.245 ;
        RECT 80.505 84.810 85.850 85.245 ;
        RECT 51.985 82.695 57.330 83.240 ;
        RECT 57.505 82.695 62.850 83.240 ;
        RECT 63.485 82.695 63.775 83.420 ;
        RECT 65.530 83.240 65.870 84.070 ;
        RECT 67.350 83.560 67.700 84.810 ;
        RECT 71.050 83.240 71.390 84.070 ;
        RECT 72.870 83.560 73.220 84.810 ;
        RECT 76.570 83.240 76.910 84.070 ;
        RECT 78.390 83.560 78.740 84.810 ;
        RECT 82.090 83.240 82.430 84.070 ;
        RECT 83.910 83.560 84.260 84.810 ;
        RECT 86.025 84.155 88.615 85.245 ;
        RECT 86.025 83.465 87.235 83.985 ;
        RECT 87.405 83.635 88.615 84.155 ;
        RECT 89.245 84.080 89.535 85.245 ;
        RECT 89.705 84.810 95.050 85.245 ;
        RECT 95.225 84.810 100.570 85.245 ;
        RECT 100.745 84.810 106.090 85.245 ;
        RECT 106.265 84.810 111.610 85.245 ;
        RECT 63.945 82.695 69.290 83.240 ;
        RECT 69.465 82.695 74.810 83.240 ;
        RECT 74.985 82.695 80.330 83.240 ;
        RECT 80.505 82.695 85.850 83.240 ;
        RECT 86.025 82.695 88.615 83.465 ;
        RECT 89.245 82.695 89.535 83.420 ;
        RECT 91.290 83.240 91.630 84.070 ;
        RECT 93.110 83.560 93.460 84.810 ;
        RECT 96.810 83.240 97.150 84.070 ;
        RECT 98.630 83.560 98.980 84.810 ;
        RECT 102.330 83.240 102.670 84.070 ;
        RECT 104.150 83.560 104.500 84.810 ;
        RECT 107.850 83.240 108.190 84.070 ;
        RECT 109.670 83.560 110.020 84.810 ;
        RECT 111.785 84.155 114.375 85.245 ;
        RECT 111.785 83.465 112.995 83.985 ;
        RECT 113.165 83.635 114.375 84.155 ;
        RECT 115.005 84.080 115.295 85.245 ;
        RECT 115.465 84.810 120.810 85.245 ;
        RECT 120.985 84.810 126.330 85.245 ;
        RECT 126.505 84.810 131.850 85.245 ;
        RECT 132.025 84.810 137.370 85.245 ;
        RECT 89.705 82.695 95.050 83.240 ;
        RECT 95.225 82.695 100.570 83.240 ;
        RECT 100.745 82.695 106.090 83.240 ;
        RECT 106.265 82.695 111.610 83.240 ;
        RECT 111.785 82.695 114.375 83.465 ;
        RECT 115.005 82.695 115.295 83.420 ;
        RECT 117.050 83.240 117.390 84.070 ;
        RECT 118.870 83.560 119.220 84.810 ;
        RECT 122.570 83.240 122.910 84.070 ;
        RECT 124.390 83.560 124.740 84.810 ;
        RECT 128.090 83.240 128.430 84.070 ;
        RECT 129.910 83.560 130.260 84.810 ;
        RECT 133.610 83.240 133.950 84.070 ;
        RECT 135.430 83.560 135.780 84.810 ;
        RECT 138.005 84.155 139.215 85.245 ;
        RECT 138.005 83.615 138.525 84.155 ;
        RECT 138.695 83.445 139.215 83.985 ;
        RECT 115.465 82.695 120.810 83.240 ;
        RECT 120.985 82.695 126.330 83.240 ;
        RECT 126.505 82.695 131.850 83.240 ;
        RECT 132.025 82.695 137.370 83.240 ;
        RECT 138.005 82.695 139.215 83.445 ;
        RECT 50.520 82.525 139.300 82.695 ;
        RECT 50.605 81.775 51.815 82.525 ;
        RECT 51.985 81.980 57.330 82.525 ;
        RECT 57.505 81.980 62.850 82.525 ;
        RECT 63.025 81.980 68.370 82.525 ;
        RECT 68.545 81.980 73.890 82.525 ;
        RECT 50.605 81.235 51.125 81.775 ;
        RECT 51.295 81.065 51.815 81.605 ;
        RECT 53.570 81.150 53.910 81.980 ;
        RECT 50.605 79.975 51.815 81.065 ;
        RECT 55.390 80.410 55.740 81.660 ;
        RECT 59.090 81.150 59.430 81.980 ;
        RECT 60.910 80.410 61.260 81.660 ;
        RECT 64.610 81.150 64.950 81.980 ;
        RECT 66.430 80.410 66.780 81.660 ;
        RECT 70.130 81.150 70.470 81.980 ;
        RECT 74.065 81.755 75.735 82.525 ;
        RECT 76.365 81.800 76.655 82.525 ;
        RECT 76.825 81.980 82.170 82.525 ;
        RECT 82.345 81.980 87.690 82.525 ;
        RECT 87.865 81.980 93.210 82.525 ;
        RECT 93.385 81.980 98.730 82.525 ;
        RECT 71.950 80.410 72.300 81.660 ;
        RECT 74.065 81.235 74.815 81.755 ;
        RECT 74.985 81.065 75.735 81.585 ;
        RECT 78.410 81.150 78.750 81.980 ;
        RECT 51.985 79.975 57.330 80.410 ;
        RECT 57.505 79.975 62.850 80.410 ;
        RECT 63.025 79.975 68.370 80.410 ;
        RECT 68.545 79.975 73.890 80.410 ;
        RECT 74.065 79.975 75.735 81.065 ;
        RECT 76.365 79.975 76.655 81.140 ;
        RECT 80.230 80.410 80.580 81.660 ;
        RECT 83.930 81.150 84.270 81.980 ;
        RECT 85.750 80.410 86.100 81.660 ;
        RECT 89.450 81.150 89.790 81.980 ;
        RECT 91.270 80.410 91.620 81.660 ;
        RECT 94.970 81.150 95.310 81.980 ;
        RECT 98.905 81.755 101.495 82.525 ;
        RECT 102.125 81.800 102.415 82.525 ;
        RECT 102.585 81.980 107.930 82.525 ;
        RECT 108.105 81.980 113.450 82.525 ;
        RECT 113.625 81.980 118.970 82.525 ;
        RECT 119.145 81.980 124.490 82.525 ;
        RECT 96.790 80.410 97.140 81.660 ;
        RECT 98.905 81.235 100.115 81.755 ;
        RECT 100.285 81.065 101.495 81.585 ;
        RECT 104.170 81.150 104.510 81.980 ;
        RECT 76.825 79.975 82.170 80.410 ;
        RECT 82.345 79.975 87.690 80.410 ;
        RECT 87.865 79.975 93.210 80.410 ;
        RECT 93.385 79.975 98.730 80.410 ;
        RECT 98.905 79.975 101.495 81.065 ;
        RECT 102.125 79.975 102.415 81.140 ;
        RECT 105.990 80.410 106.340 81.660 ;
        RECT 109.690 81.150 110.030 81.980 ;
        RECT 111.510 80.410 111.860 81.660 ;
        RECT 115.210 81.150 115.550 81.980 ;
        RECT 117.030 80.410 117.380 81.660 ;
        RECT 120.730 81.150 121.070 81.980 ;
        RECT 124.665 81.755 127.255 82.525 ;
        RECT 127.885 81.800 128.175 82.525 ;
        RECT 128.345 81.980 133.690 82.525 ;
        RECT 122.550 80.410 122.900 81.660 ;
        RECT 124.665 81.235 125.875 81.755 ;
        RECT 126.045 81.065 127.255 81.585 ;
        RECT 129.930 81.150 130.270 81.980 ;
        RECT 133.865 81.755 137.375 82.525 ;
        RECT 138.005 81.775 139.215 82.525 ;
        RECT 102.585 79.975 107.930 80.410 ;
        RECT 108.105 79.975 113.450 80.410 ;
        RECT 113.625 79.975 118.970 80.410 ;
        RECT 119.145 79.975 124.490 80.410 ;
        RECT 124.665 79.975 127.255 81.065 ;
        RECT 127.885 79.975 128.175 81.140 ;
        RECT 131.750 80.410 132.100 81.660 ;
        RECT 133.865 81.235 135.515 81.755 ;
        RECT 135.685 81.065 137.375 81.585 ;
        RECT 128.345 79.975 133.690 80.410 ;
        RECT 133.865 79.975 137.375 81.065 ;
        RECT 138.005 81.065 138.525 81.605 ;
        RECT 138.695 81.235 139.215 81.775 ;
        RECT 138.005 79.975 139.215 81.065 ;
        RECT 50.520 79.805 139.300 79.975 ;
        RECT 50.605 78.715 51.815 79.805 ;
        RECT 51.985 79.370 57.330 79.805 ;
        RECT 57.505 79.370 62.850 79.805 ;
        RECT 50.605 78.005 51.125 78.545 ;
        RECT 51.295 78.175 51.815 78.715 ;
        RECT 50.605 77.255 51.815 78.005 ;
        RECT 53.570 77.800 53.910 78.630 ;
        RECT 55.390 78.120 55.740 79.370 ;
        RECT 59.090 77.800 59.430 78.630 ;
        RECT 60.910 78.120 61.260 79.370 ;
        RECT 63.485 78.640 63.775 79.805 ;
        RECT 63.945 79.370 69.290 79.805 ;
        RECT 69.465 79.370 74.810 79.805 ;
        RECT 74.985 79.370 80.330 79.805 ;
        RECT 80.505 79.370 85.850 79.805 ;
        RECT 51.985 77.255 57.330 77.800 ;
        RECT 57.505 77.255 62.850 77.800 ;
        RECT 63.485 77.255 63.775 77.980 ;
        RECT 65.530 77.800 65.870 78.630 ;
        RECT 67.350 78.120 67.700 79.370 ;
        RECT 71.050 77.800 71.390 78.630 ;
        RECT 72.870 78.120 73.220 79.370 ;
        RECT 76.570 77.800 76.910 78.630 ;
        RECT 78.390 78.120 78.740 79.370 ;
        RECT 82.090 77.800 82.430 78.630 ;
        RECT 83.910 78.120 84.260 79.370 ;
        RECT 86.025 78.715 88.615 79.805 ;
        RECT 86.025 78.025 87.235 78.545 ;
        RECT 87.405 78.195 88.615 78.715 ;
        RECT 89.245 78.640 89.535 79.805 ;
        RECT 89.705 79.370 95.050 79.805 ;
        RECT 95.225 79.370 100.570 79.805 ;
        RECT 100.745 79.370 106.090 79.805 ;
        RECT 106.265 79.370 111.610 79.805 ;
        RECT 63.945 77.255 69.290 77.800 ;
        RECT 69.465 77.255 74.810 77.800 ;
        RECT 74.985 77.255 80.330 77.800 ;
        RECT 80.505 77.255 85.850 77.800 ;
        RECT 86.025 77.255 88.615 78.025 ;
        RECT 89.245 77.255 89.535 77.980 ;
        RECT 91.290 77.800 91.630 78.630 ;
        RECT 93.110 78.120 93.460 79.370 ;
        RECT 96.810 77.800 97.150 78.630 ;
        RECT 98.630 78.120 98.980 79.370 ;
        RECT 102.330 77.800 102.670 78.630 ;
        RECT 104.150 78.120 104.500 79.370 ;
        RECT 107.850 77.800 108.190 78.630 ;
        RECT 109.670 78.120 110.020 79.370 ;
        RECT 111.785 78.715 114.375 79.805 ;
        RECT 111.785 78.025 112.995 78.545 ;
        RECT 113.165 78.195 114.375 78.715 ;
        RECT 115.005 78.640 115.295 79.805 ;
        RECT 115.465 79.370 120.810 79.805 ;
        RECT 120.985 79.370 126.330 79.805 ;
        RECT 126.505 79.370 131.850 79.805 ;
        RECT 132.025 79.370 137.370 79.805 ;
        RECT 89.705 77.255 95.050 77.800 ;
        RECT 95.225 77.255 100.570 77.800 ;
        RECT 100.745 77.255 106.090 77.800 ;
        RECT 106.265 77.255 111.610 77.800 ;
        RECT 111.785 77.255 114.375 78.025 ;
        RECT 115.005 77.255 115.295 77.980 ;
        RECT 117.050 77.800 117.390 78.630 ;
        RECT 118.870 78.120 119.220 79.370 ;
        RECT 122.570 77.800 122.910 78.630 ;
        RECT 124.390 78.120 124.740 79.370 ;
        RECT 128.090 77.800 128.430 78.630 ;
        RECT 129.910 78.120 130.260 79.370 ;
        RECT 133.610 77.800 133.950 78.630 ;
        RECT 135.430 78.120 135.780 79.370 ;
        RECT 138.005 78.715 139.215 79.805 ;
        RECT 138.005 78.175 138.525 78.715 ;
        RECT 138.695 78.005 139.215 78.545 ;
        RECT 115.465 77.255 120.810 77.800 ;
        RECT 120.985 77.255 126.330 77.800 ;
        RECT 126.505 77.255 131.850 77.800 ;
        RECT 132.025 77.255 137.370 77.800 ;
        RECT 138.005 77.255 139.215 78.005 ;
        RECT 50.520 77.085 139.300 77.255 ;
        RECT 50.605 76.335 51.815 77.085 ;
        RECT 51.985 76.540 57.330 77.085 ;
        RECT 57.505 76.540 62.850 77.085 ;
        RECT 63.025 76.540 68.370 77.085 ;
        RECT 68.545 76.540 73.890 77.085 ;
        RECT 50.605 75.795 51.125 76.335 ;
        RECT 51.295 75.625 51.815 76.165 ;
        RECT 53.570 75.710 53.910 76.540 ;
        RECT 50.605 74.535 51.815 75.625 ;
        RECT 55.390 74.970 55.740 76.220 ;
        RECT 59.090 75.710 59.430 76.540 ;
        RECT 60.910 74.970 61.260 76.220 ;
        RECT 64.610 75.710 64.950 76.540 ;
        RECT 66.430 74.970 66.780 76.220 ;
        RECT 70.130 75.710 70.470 76.540 ;
        RECT 74.065 76.315 75.735 77.085 ;
        RECT 76.365 76.360 76.655 77.085 ;
        RECT 76.825 76.540 82.170 77.085 ;
        RECT 82.345 76.540 87.690 77.085 ;
        RECT 87.865 76.540 93.210 77.085 ;
        RECT 93.385 76.540 98.730 77.085 ;
        RECT 71.950 74.970 72.300 76.220 ;
        RECT 74.065 75.795 74.815 76.315 ;
        RECT 74.985 75.625 75.735 76.145 ;
        RECT 78.410 75.710 78.750 76.540 ;
        RECT 51.985 74.535 57.330 74.970 ;
        RECT 57.505 74.535 62.850 74.970 ;
        RECT 63.025 74.535 68.370 74.970 ;
        RECT 68.545 74.535 73.890 74.970 ;
        RECT 74.065 74.535 75.735 75.625 ;
        RECT 76.365 74.535 76.655 75.700 ;
        RECT 80.230 74.970 80.580 76.220 ;
        RECT 83.930 75.710 84.270 76.540 ;
        RECT 85.750 74.970 86.100 76.220 ;
        RECT 89.450 75.710 89.790 76.540 ;
        RECT 91.270 74.970 91.620 76.220 ;
        RECT 94.970 75.710 95.310 76.540 ;
        RECT 98.905 76.315 101.495 77.085 ;
        RECT 102.125 76.360 102.415 77.085 ;
        RECT 102.585 76.540 107.930 77.085 ;
        RECT 108.105 76.540 113.450 77.085 ;
        RECT 113.625 76.540 118.970 77.085 ;
        RECT 119.145 76.540 124.490 77.085 ;
        RECT 96.790 74.970 97.140 76.220 ;
        RECT 98.905 75.795 100.115 76.315 ;
        RECT 100.285 75.625 101.495 76.145 ;
        RECT 104.170 75.710 104.510 76.540 ;
        RECT 76.825 74.535 82.170 74.970 ;
        RECT 82.345 74.535 87.690 74.970 ;
        RECT 87.865 74.535 93.210 74.970 ;
        RECT 93.385 74.535 98.730 74.970 ;
        RECT 98.905 74.535 101.495 75.625 ;
        RECT 102.125 74.535 102.415 75.700 ;
        RECT 105.990 74.970 106.340 76.220 ;
        RECT 109.690 75.710 110.030 76.540 ;
        RECT 111.510 74.970 111.860 76.220 ;
        RECT 115.210 75.710 115.550 76.540 ;
        RECT 117.030 74.970 117.380 76.220 ;
        RECT 120.730 75.710 121.070 76.540 ;
        RECT 124.665 76.315 127.255 77.085 ;
        RECT 127.885 76.360 128.175 77.085 ;
        RECT 128.345 76.540 133.690 77.085 ;
        RECT 122.550 74.970 122.900 76.220 ;
        RECT 124.665 75.795 125.875 76.315 ;
        RECT 126.045 75.625 127.255 76.145 ;
        RECT 129.930 75.710 130.270 76.540 ;
        RECT 133.865 76.315 137.375 77.085 ;
        RECT 138.005 76.335 139.215 77.085 ;
        RECT 102.585 74.535 107.930 74.970 ;
        RECT 108.105 74.535 113.450 74.970 ;
        RECT 113.625 74.535 118.970 74.970 ;
        RECT 119.145 74.535 124.490 74.970 ;
        RECT 124.665 74.535 127.255 75.625 ;
        RECT 127.885 74.535 128.175 75.700 ;
        RECT 131.750 74.970 132.100 76.220 ;
        RECT 133.865 75.795 135.515 76.315 ;
        RECT 135.685 75.625 137.375 76.145 ;
        RECT 128.345 74.535 133.690 74.970 ;
        RECT 133.865 74.535 137.375 75.625 ;
        RECT 138.005 75.625 138.525 76.165 ;
        RECT 138.695 75.795 139.215 76.335 ;
        RECT 138.005 74.535 139.215 75.625 ;
        RECT 50.520 74.365 139.300 74.535 ;
        RECT 50.605 73.275 51.815 74.365 ;
        RECT 51.985 73.930 57.330 74.365 ;
        RECT 57.505 73.930 62.850 74.365 ;
        RECT 50.605 72.565 51.125 73.105 ;
        RECT 51.295 72.735 51.815 73.275 ;
        RECT 50.605 71.815 51.815 72.565 ;
        RECT 53.570 72.360 53.910 73.190 ;
        RECT 55.390 72.680 55.740 73.930 ;
        RECT 59.090 72.360 59.430 73.190 ;
        RECT 60.910 72.680 61.260 73.930 ;
        RECT 63.485 73.200 63.775 74.365 ;
        RECT 63.945 73.930 69.290 74.365 ;
        RECT 69.465 73.930 74.810 74.365 ;
        RECT 74.985 73.930 80.330 74.365 ;
        RECT 80.505 73.930 85.850 74.365 ;
        RECT 51.985 71.815 57.330 72.360 ;
        RECT 57.505 71.815 62.850 72.360 ;
        RECT 63.485 71.815 63.775 72.540 ;
        RECT 65.530 72.360 65.870 73.190 ;
        RECT 67.350 72.680 67.700 73.930 ;
        RECT 71.050 72.360 71.390 73.190 ;
        RECT 72.870 72.680 73.220 73.930 ;
        RECT 76.570 72.360 76.910 73.190 ;
        RECT 78.390 72.680 78.740 73.930 ;
        RECT 82.090 72.360 82.430 73.190 ;
        RECT 83.910 72.680 84.260 73.930 ;
        RECT 86.025 73.275 88.615 74.365 ;
        RECT 86.025 72.585 87.235 73.105 ;
        RECT 87.405 72.755 88.615 73.275 ;
        RECT 89.245 73.200 89.535 74.365 ;
        RECT 89.705 73.930 95.050 74.365 ;
        RECT 95.225 73.930 100.570 74.365 ;
        RECT 100.745 73.930 106.090 74.365 ;
        RECT 106.265 73.930 111.610 74.365 ;
        RECT 63.945 71.815 69.290 72.360 ;
        RECT 69.465 71.815 74.810 72.360 ;
        RECT 74.985 71.815 80.330 72.360 ;
        RECT 80.505 71.815 85.850 72.360 ;
        RECT 86.025 71.815 88.615 72.585 ;
        RECT 89.245 71.815 89.535 72.540 ;
        RECT 91.290 72.360 91.630 73.190 ;
        RECT 93.110 72.680 93.460 73.930 ;
        RECT 96.810 72.360 97.150 73.190 ;
        RECT 98.630 72.680 98.980 73.930 ;
        RECT 102.330 72.360 102.670 73.190 ;
        RECT 104.150 72.680 104.500 73.930 ;
        RECT 107.850 72.360 108.190 73.190 ;
        RECT 109.670 72.680 110.020 73.930 ;
        RECT 111.785 73.275 114.375 74.365 ;
        RECT 111.785 72.585 112.995 73.105 ;
        RECT 113.165 72.755 114.375 73.275 ;
        RECT 115.005 73.200 115.295 74.365 ;
        RECT 115.465 73.930 120.810 74.365 ;
        RECT 120.985 73.930 126.330 74.365 ;
        RECT 126.505 73.930 131.850 74.365 ;
        RECT 132.025 73.930 137.370 74.365 ;
        RECT 89.705 71.815 95.050 72.360 ;
        RECT 95.225 71.815 100.570 72.360 ;
        RECT 100.745 71.815 106.090 72.360 ;
        RECT 106.265 71.815 111.610 72.360 ;
        RECT 111.785 71.815 114.375 72.585 ;
        RECT 115.005 71.815 115.295 72.540 ;
        RECT 117.050 72.360 117.390 73.190 ;
        RECT 118.870 72.680 119.220 73.930 ;
        RECT 122.570 72.360 122.910 73.190 ;
        RECT 124.390 72.680 124.740 73.930 ;
        RECT 128.090 72.360 128.430 73.190 ;
        RECT 129.910 72.680 130.260 73.930 ;
        RECT 133.610 72.360 133.950 73.190 ;
        RECT 135.430 72.680 135.780 73.930 ;
        RECT 138.005 73.275 139.215 74.365 ;
        RECT 138.005 72.735 138.525 73.275 ;
        RECT 138.695 72.565 139.215 73.105 ;
        RECT 115.465 71.815 120.810 72.360 ;
        RECT 120.985 71.815 126.330 72.360 ;
        RECT 126.505 71.815 131.850 72.360 ;
        RECT 132.025 71.815 137.370 72.360 ;
        RECT 138.005 71.815 139.215 72.565 ;
        RECT 50.520 71.645 139.300 71.815 ;
        RECT 50.605 70.895 51.815 71.645 ;
        RECT 51.985 71.100 57.330 71.645 ;
        RECT 57.505 71.100 62.850 71.645 ;
        RECT 63.025 71.100 68.370 71.645 ;
        RECT 68.545 71.100 73.890 71.645 ;
        RECT 50.605 70.355 51.125 70.895 ;
        RECT 51.295 70.185 51.815 70.725 ;
        RECT 53.570 70.270 53.910 71.100 ;
        RECT 50.605 69.095 51.815 70.185 ;
        RECT 55.390 69.530 55.740 70.780 ;
        RECT 59.090 70.270 59.430 71.100 ;
        RECT 60.910 69.530 61.260 70.780 ;
        RECT 64.610 70.270 64.950 71.100 ;
        RECT 66.430 69.530 66.780 70.780 ;
        RECT 70.130 70.270 70.470 71.100 ;
        RECT 74.065 70.875 75.735 71.645 ;
        RECT 76.365 70.920 76.655 71.645 ;
        RECT 76.825 71.100 82.170 71.645 ;
        RECT 82.345 71.100 87.690 71.645 ;
        RECT 87.865 71.100 93.210 71.645 ;
        RECT 93.385 71.100 98.730 71.645 ;
        RECT 71.950 69.530 72.300 70.780 ;
        RECT 74.065 70.355 74.815 70.875 ;
        RECT 74.985 70.185 75.735 70.705 ;
        RECT 78.410 70.270 78.750 71.100 ;
        RECT 51.985 69.095 57.330 69.530 ;
        RECT 57.505 69.095 62.850 69.530 ;
        RECT 63.025 69.095 68.370 69.530 ;
        RECT 68.545 69.095 73.890 69.530 ;
        RECT 74.065 69.095 75.735 70.185 ;
        RECT 76.365 69.095 76.655 70.260 ;
        RECT 80.230 69.530 80.580 70.780 ;
        RECT 83.930 70.270 84.270 71.100 ;
        RECT 85.750 69.530 86.100 70.780 ;
        RECT 89.450 70.270 89.790 71.100 ;
        RECT 91.270 69.530 91.620 70.780 ;
        RECT 94.970 70.270 95.310 71.100 ;
        RECT 98.905 70.875 101.495 71.645 ;
        RECT 102.125 70.920 102.415 71.645 ;
        RECT 102.585 71.100 107.930 71.645 ;
        RECT 108.105 71.100 113.450 71.645 ;
        RECT 113.625 71.100 118.970 71.645 ;
        RECT 119.145 71.100 124.490 71.645 ;
        RECT 96.790 69.530 97.140 70.780 ;
        RECT 98.905 70.355 100.115 70.875 ;
        RECT 100.285 70.185 101.495 70.705 ;
        RECT 104.170 70.270 104.510 71.100 ;
        RECT 76.825 69.095 82.170 69.530 ;
        RECT 82.345 69.095 87.690 69.530 ;
        RECT 87.865 69.095 93.210 69.530 ;
        RECT 93.385 69.095 98.730 69.530 ;
        RECT 98.905 69.095 101.495 70.185 ;
        RECT 102.125 69.095 102.415 70.260 ;
        RECT 105.990 69.530 106.340 70.780 ;
        RECT 109.690 70.270 110.030 71.100 ;
        RECT 111.510 69.530 111.860 70.780 ;
        RECT 115.210 70.270 115.550 71.100 ;
        RECT 117.030 69.530 117.380 70.780 ;
        RECT 120.730 70.270 121.070 71.100 ;
        RECT 124.665 70.875 127.255 71.645 ;
        RECT 127.885 70.920 128.175 71.645 ;
        RECT 128.345 71.100 133.690 71.645 ;
        RECT 122.550 69.530 122.900 70.780 ;
        RECT 124.665 70.355 125.875 70.875 ;
        RECT 126.045 70.185 127.255 70.705 ;
        RECT 129.930 70.270 130.270 71.100 ;
        RECT 133.865 70.875 137.375 71.645 ;
        RECT 138.005 70.895 139.215 71.645 ;
        RECT 102.585 69.095 107.930 69.530 ;
        RECT 108.105 69.095 113.450 69.530 ;
        RECT 113.625 69.095 118.970 69.530 ;
        RECT 119.145 69.095 124.490 69.530 ;
        RECT 124.665 69.095 127.255 70.185 ;
        RECT 127.885 69.095 128.175 70.260 ;
        RECT 131.750 69.530 132.100 70.780 ;
        RECT 133.865 70.355 135.515 70.875 ;
        RECT 135.685 70.185 137.375 70.705 ;
        RECT 128.345 69.095 133.690 69.530 ;
        RECT 133.865 69.095 137.375 70.185 ;
        RECT 138.005 70.185 138.525 70.725 ;
        RECT 138.695 70.355 139.215 70.895 ;
        RECT 138.005 69.095 139.215 70.185 ;
        RECT 50.520 68.925 139.300 69.095 ;
        RECT 50.605 67.835 51.815 68.925 ;
        RECT 51.985 68.490 57.330 68.925 ;
        RECT 57.505 68.490 62.850 68.925 ;
        RECT 50.605 67.125 51.125 67.665 ;
        RECT 51.295 67.295 51.815 67.835 ;
        RECT 50.605 66.375 51.815 67.125 ;
        RECT 53.570 66.920 53.910 67.750 ;
        RECT 55.390 67.240 55.740 68.490 ;
        RECT 59.090 66.920 59.430 67.750 ;
        RECT 60.910 67.240 61.260 68.490 ;
        RECT 63.485 67.760 63.775 68.925 ;
        RECT 63.945 68.490 69.290 68.925 ;
        RECT 69.465 68.490 74.810 68.925 ;
        RECT 74.985 68.490 80.330 68.925 ;
        RECT 80.505 68.490 85.850 68.925 ;
        RECT 51.985 66.375 57.330 66.920 ;
        RECT 57.505 66.375 62.850 66.920 ;
        RECT 63.485 66.375 63.775 67.100 ;
        RECT 65.530 66.920 65.870 67.750 ;
        RECT 67.350 67.240 67.700 68.490 ;
        RECT 71.050 66.920 71.390 67.750 ;
        RECT 72.870 67.240 73.220 68.490 ;
        RECT 76.570 66.920 76.910 67.750 ;
        RECT 78.390 67.240 78.740 68.490 ;
        RECT 82.090 66.920 82.430 67.750 ;
        RECT 83.910 67.240 84.260 68.490 ;
        RECT 86.025 67.835 88.615 68.925 ;
        RECT 86.025 67.145 87.235 67.665 ;
        RECT 87.405 67.315 88.615 67.835 ;
        RECT 89.245 67.760 89.535 68.925 ;
        RECT 89.705 68.490 95.050 68.925 ;
        RECT 95.225 68.490 100.570 68.925 ;
        RECT 100.745 68.490 106.090 68.925 ;
        RECT 106.265 68.490 111.610 68.925 ;
        RECT 63.945 66.375 69.290 66.920 ;
        RECT 69.465 66.375 74.810 66.920 ;
        RECT 74.985 66.375 80.330 66.920 ;
        RECT 80.505 66.375 85.850 66.920 ;
        RECT 86.025 66.375 88.615 67.145 ;
        RECT 89.245 66.375 89.535 67.100 ;
        RECT 91.290 66.920 91.630 67.750 ;
        RECT 93.110 67.240 93.460 68.490 ;
        RECT 96.810 66.920 97.150 67.750 ;
        RECT 98.630 67.240 98.980 68.490 ;
        RECT 102.330 66.920 102.670 67.750 ;
        RECT 104.150 67.240 104.500 68.490 ;
        RECT 107.850 66.920 108.190 67.750 ;
        RECT 109.670 67.240 110.020 68.490 ;
        RECT 111.785 67.835 114.375 68.925 ;
        RECT 111.785 67.145 112.995 67.665 ;
        RECT 113.165 67.315 114.375 67.835 ;
        RECT 115.005 67.760 115.295 68.925 ;
        RECT 115.465 68.490 120.810 68.925 ;
        RECT 120.985 68.490 126.330 68.925 ;
        RECT 126.505 68.490 131.850 68.925 ;
        RECT 132.025 68.490 137.370 68.925 ;
        RECT 89.705 66.375 95.050 66.920 ;
        RECT 95.225 66.375 100.570 66.920 ;
        RECT 100.745 66.375 106.090 66.920 ;
        RECT 106.265 66.375 111.610 66.920 ;
        RECT 111.785 66.375 114.375 67.145 ;
        RECT 115.005 66.375 115.295 67.100 ;
        RECT 117.050 66.920 117.390 67.750 ;
        RECT 118.870 67.240 119.220 68.490 ;
        RECT 122.570 66.920 122.910 67.750 ;
        RECT 124.390 67.240 124.740 68.490 ;
        RECT 128.090 66.920 128.430 67.750 ;
        RECT 129.910 67.240 130.260 68.490 ;
        RECT 133.610 66.920 133.950 67.750 ;
        RECT 135.430 67.240 135.780 68.490 ;
        RECT 138.005 67.835 139.215 68.925 ;
        RECT 138.005 67.295 138.525 67.835 ;
        RECT 138.695 67.125 139.215 67.665 ;
        RECT 115.465 66.375 120.810 66.920 ;
        RECT 120.985 66.375 126.330 66.920 ;
        RECT 126.505 66.375 131.850 66.920 ;
        RECT 132.025 66.375 137.370 66.920 ;
        RECT 138.005 66.375 139.215 67.125 ;
        RECT 50.520 66.205 139.300 66.375 ;
        RECT 50.605 65.455 51.815 66.205 ;
        RECT 51.985 65.660 57.330 66.205 ;
        RECT 57.505 65.660 62.850 66.205 ;
        RECT 63.025 65.660 68.370 66.205 ;
        RECT 68.545 65.660 73.890 66.205 ;
        RECT 50.605 64.915 51.125 65.455 ;
        RECT 51.295 64.745 51.815 65.285 ;
        RECT 53.570 64.830 53.910 65.660 ;
        RECT 50.605 63.655 51.815 64.745 ;
        RECT 55.390 64.090 55.740 65.340 ;
        RECT 59.090 64.830 59.430 65.660 ;
        RECT 60.910 64.090 61.260 65.340 ;
        RECT 64.610 64.830 64.950 65.660 ;
        RECT 66.430 64.090 66.780 65.340 ;
        RECT 70.130 64.830 70.470 65.660 ;
        RECT 74.065 65.435 75.735 66.205 ;
        RECT 76.365 65.480 76.655 66.205 ;
        RECT 76.825 65.660 82.170 66.205 ;
        RECT 82.345 65.660 87.690 66.205 ;
        RECT 87.865 65.660 93.210 66.205 ;
        RECT 93.385 65.660 98.730 66.205 ;
        RECT 71.950 64.090 72.300 65.340 ;
        RECT 74.065 64.915 74.815 65.435 ;
        RECT 74.985 64.745 75.735 65.265 ;
        RECT 78.410 64.830 78.750 65.660 ;
        RECT 51.985 63.655 57.330 64.090 ;
        RECT 57.505 63.655 62.850 64.090 ;
        RECT 63.025 63.655 68.370 64.090 ;
        RECT 68.545 63.655 73.890 64.090 ;
        RECT 74.065 63.655 75.735 64.745 ;
        RECT 76.365 63.655 76.655 64.820 ;
        RECT 80.230 64.090 80.580 65.340 ;
        RECT 83.930 64.830 84.270 65.660 ;
        RECT 85.750 64.090 86.100 65.340 ;
        RECT 89.450 64.830 89.790 65.660 ;
        RECT 91.270 64.090 91.620 65.340 ;
        RECT 94.970 64.830 95.310 65.660 ;
        RECT 98.905 65.435 101.495 66.205 ;
        RECT 102.125 65.480 102.415 66.205 ;
        RECT 102.585 65.660 107.930 66.205 ;
        RECT 108.105 65.660 113.450 66.205 ;
        RECT 113.625 65.660 118.970 66.205 ;
        RECT 119.145 65.660 124.490 66.205 ;
        RECT 96.790 64.090 97.140 65.340 ;
        RECT 98.905 64.915 100.115 65.435 ;
        RECT 100.285 64.745 101.495 65.265 ;
        RECT 104.170 64.830 104.510 65.660 ;
        RECT 76.825 63.655 82.170 64.090 ;
        RECT 82.345 63.655 87.690 64.090 ;
        RECT 87.865 63.655 93.210 64.090 ;
        RECT 93.385 63.655 98.730 64.090 ;
        RECT 98.905 63.655 101.495 64.745 ;
        RECT 102.125 63.655 102.415 64.820 ;
        RECT 105.990 64.090 106.340 65.340 ;
        RECT 109.690 64.830 110.030 65.660 ;
        RECT 111.510 64.090 111.860 65.340 ;
        RECT 115.210 64.830 115.550 65.660 ;
        RECT 117.030 64.090 117.380 65.340 ;
        RECT 120.730 64.830 121.070 65.660 ;
        RECT 124.665 65.435 127.255 66.205 ;
        RECT 127.885 65.480 128.175 66.205 ;
        RECT 128.345 65.660 133.690 66.205 ;
        RECT 122.550 64.090 122.900 65.340 ;
        RECT 124.665 64.915 125.875 65.435 ;
        RECT 126.045 64.745 127.255 65.265 ;
        RECT 129.930 64.830 130.270 65.660 ;
        RECT 133.865 65.435 137.375 66.205 ;
        RECT 138.005 65.455 139.215 66.205 ;
        RECT 102.585 63.655 107.930 64.090 ;
        RECT 108.105 63.655 113.450 64.090 ;
        RECT 113.625 63.655 118.970 64.090 ;
        RECT 119.145 63.655 124.490 64.090 ;
        RECT 124.665 63.655 127.255 64.745 ;
        RECT 127.885 63.655 128.175 64.820 ;
        RECT 131.750 64.090 132.100 65.340 ;
        RECT 133.865 64.915 135.515 65.435 ;
        RECT 135.685 64.745 137.375 65.265 ;
        RECT 128.345 63.655 133.690 64.090 ;
        RECT 133.865 63.655 137.375 64.745 ;
        RECT 138.005 64.745 138.525 65.285 ;
        RECT 138.695 64.915 139.215 65.455 ;
        RECT 138.005 63.655 139.215 64.745 ;
        RECT 50.520 63.485 139.300 63.655 ;
        RECT 50.605 62.395 51.815 63.485 ;
        RECT 51.985 63.050 57.330 63.485 ;
        RECT 57.505 63.050 62.850 63.485 ;
        RECT 50.605 61.685 51.125 62.225 ;
        RECT 51.295 61.855 51.815 62.395 ;
        RECT 50.605 60.935 51.815 61.685 ;
        RECT 53.570 61.480 53.910 62.310 ;
        RECT 55.390 61.800 55.740 63.050 ;
        RECT 59.090 61.480 59.430 62.310 ;
        RECT 60.910 61.800 61.260 63.050 ;
        RECT 63.485 62.320 63.775 63.485 ;
        RECT 63.945 63.050 69.290 63.485 ;
        RECT 69.465 63.050 74.810 63.485 ;
        RECT 51.985 60.935 57.330 61.480 ;
        RECT 57.505 60.935 62.850 61.480 ;
        RECT 63.485 60.935 63.775 61.660 ;
        RECT 65.530 61.480 65.870 62.310 ;
        RECT 67.350 61.800 67.700 63.050 ;
        RECT 71.050 61.480 71.390 62.310 ;
        RECT 72.870 61.800 73.220 63.050 ;
        RECT 74.985 62.395 76.195 63.485 ;
        RECT 74.985 61.685 75.505 62.225 ;
        RECT 75.675 61.855 76.195 62.395 ;
        RECT 76.365 62.320 76.655 63.485 ;
        RECT 76.825 63.050 82.170 63.485 ;
        RECT 82.345 63.050 87.690 63.485 ;
        RECT 63.945 60.935 69.290 61.480 ;
        RECT 69.465 60.935 74.810 61.480 ;
        RECT 74.985 60.935 76.195 61.685 ;
        RECT 76.365 60.935 76.655 61.660 ;
        RECT 78.410 61.480 78.750 62.310 ;
        RECT 80.230 61.800 80.580 63.050 ;
        RECT 83.930 61.480 84.270 62.310 ;
        RECT 85.750 61.800 86.100 63.050 ;
        RECT 87.865 62.395 89.075 63.485 ;
        RECT 87.865 61.685 88.385 62.225 ;
        RECT 88.555 61.855 89.075 62.395 ;
        RECT 89.245 62.320 89.535 63.485 ;
        RECT 89.705 63.050 95.050 63.485 ;
        RECT 95.225 63.050 100.570 63.485 ;
        RECT 76.825 60.935 82.170 61.480 ;
        RECT 82.345 60.935 87.690 61.480 ;
        RECT 87.865 60.935 89.075 61.685 ;
        RECT 89.245 60.935 89.535 61.660 ;
        RECT 91.290 61.480 91.630 62.310 ;
        RECT 93.110 61.800 93.460 63.050 ;
        RECT 96.810 61.480 97.150 62.310 ;
        RECT 98.630 61.800 98.980 63.050 ;
        RECT 100.745 62.395 101.955 63.485 ;
        RECT 100.745 61.685 101.265 62.225 ;
        RECT 101.435 61.855 101.955 62.395 ;
        RECT 102.125 62.320 102.415 63.485 ;
        RECT 102.585 63.050 107.930 63.485 ;
        RECT 108.105 63.050 113.450 63.485 ;
        RECT 89.705 60.935 95.050 61.480 ;
        RECT 95.225 60.935 100.570 61.480 ;
        RECT 100.745 60.935 101.955 61.685 ;
        RECT 102.125 60.935 102.415 61.660 ;
        RECT 104.170 61.480 104.510 62.310 ;
        RECT 105.990 61.800 106.340 63.050 ;
        RECT 109.690 61.480 110.030 62.310 ;
        RECT 111.510 61.800 111.860 63.050 ;
        RECT 113.625 62.395 114.835 63.485 ;
        RECT 113.625 61.685 114.145 62.225 ;
        RECT 114.315 61.855 114.835 62.395 ;
        RECT 115.005 62.320 115.295 63.485 ;
        RECT 115.465 63.050 120.810 63.485 ;
        RECT 120.985 63.050 126.330 63.485 ;
        RECT 102.585 60.935 107.930 61.480 ;
        RECT 108.105 60.935 113.450 61.480 ;
        RECT 113.625 60.935 114.835 61.685 ;
        RECT 115.005 60.935 115.295 61.660 ;
        RECT 117.050 61.480 117.390 62.310 ;
        RECT 118.870 61.800 119.220 63.050 ;
        RECT 122.570 61.480 122.910 62.310 ;
        RECT 124.390 61.800 124.740 63.050 ;
        RECT 126.505 62.395 127.715 63.485 ;
        RECT 126.505 61.685 127.025 62.225 ;
        RECT 127.195 61.855 127.715 62.395 ;
        RECT 127.885 62.320 128.175 63.485 ;
        RECT 128.345 63.050 133.690 63.485 ;
        RECT 115.465 60.935 120.810 61.480 ;
        RECT 120.985 60.935 126.330 61.480 ;
        RECT 126.505 60.935 127.715 61.685 ;
        RECT 127.885 60.935 128.175 61.660 ;
        RECT 129.930 61.480 130.270 62.310 ;
        RECT 131.750 61.800 132.100 63.050 ;
        RECT 133.865 62.395 137.375 63.485 ;
        RECT 133.865 61.705 135.515 62.225 ;
        RECT 135.685 61.875 137.375 62.395 ;
        RECT 138.005 62.395 139.215 63.485 ;
        RECT 138.005 61.855 138.525 62.395 ;
        RECT 128.345 60.935 133.690 61.480 ;
        RECT 133.865 60.935 137.375 61.705 ;
        RECT 138.695 61.685 139.215 62.225 ;
        RECT 138.005 60.935 139.215 61.685 ;
        RECT 50.520 60.765 139.300 60.935 ;
      LAYER mcon ;
        RECT 50.665 136.925 50.835 137.095 ;
        RECT 51.125 136.925 51.295 137.095 ;
        RECT 51.585 136.925 51.755 137.095 ;
        RECT 52.045 136.925 52.215 137.095 ;
        RECT 52.505 136.925 52.675 137.095 ;
        RECT 52.965 136.925 53.135 137.095 ;
        RECT 53.425 136.925 53.595 137.095 ;
        RECT 53.885 136.925 54.055 137.095 ;
        RECT 54.345 136.925 54.515 137.095 ;
        RECT 54.805 136.925 54.975 137.095 ;
        RECT 55.265 136.925 55.435 137.095 ;
        RECT 55.725 136.925 55.895 137.095 ;
        RECT 56.185 136.925 56.355 137.095 ;
        RECT 56.645 136.925 56.815 137.095 ;
        RECT 57.105 136.925 57.275 137.095 ;
        RECT 57.565 136.925 57.735 137.095 ;
        RECT 58.025 136.925 58.195 137.095 ;
        RECT 58.485 136.925 58.655 137.095 ;
        RECT 58.945 136.925 59.115 137.095 ;
        RECT 59.405 136.925 59.575 137.095 ;
        RECT 59.865 136.925 60.035 137.095 ;
        RECT 60.325 136.925 60.495 137.095 ;
        RECT 60.785 136.925 60.955 137.095 ;
        RECT 61.245 136.925 61.415 137.095 ;
        RECT 61.705 136.925 61.875 137.095 ;
        RECT 62.165 136.925 62.335 137.095 ;
        RECT 62.625 136.925 62.795 137.095 ;
        RECT 63.085 136.925 63.255 137.095 ;
        RECT 63.545 136.925 63.715 137.095 ;
        RECT 64.005 136.925 64.175 137.095 ;
        RECT 64.465 136.925 64.635 137.095 ;
        RECT 64.925 136.925 65.095 137.095 ;
        RECT 65.385 136.925 65.555 137.095 ;
        RECT 65.845 136.925 66.015 137.095 ;
        RECT 66.305 136.925 66.475 137.095 ;
        RECT 66.765 136.925 66.935 137.095 ;
        RECT 67.225 136.925 67.395 137.095 ;
        RECT 67.685 136.925 67.855 137.095 ;
        RECT 68.145 136.925 68.315 137.095 ;
        RECT 68.605 136.925 68.775 137.095 ;
        RECT 69.065 136.925 69.235 137.095 ;
        RECT 69.525 136.925 69.695 137.095 ;
        RECT 69.985 136.925 70.155 137.095 ;
        RECT 70.445 136.925 70.615 137.095 ;
        RECT 70.905 136.925 71.075 137.095 ;
        RECT 71.365 136.925 71.535 137.095 ;
        RECT 71.825 136.925 71.995 137.095 ;
        RECT 72.285 136.925 72.455 137.095 ;
        RECT 72.745 136.925 72.915 137.095 ;
        RECT 73.205 136.925 73.375 137.095 ;
        RECT 73.665 136.925 73.835 137.095 ;
        RECT 74.125 136.925 74.295 137.095 ;
        RECT 74.585 136.925 74.755 137.095 ;
        RECT 75.045 136.925 75.215 137.095 ;
        RECT 75.505 136.925 75.675 137.095 ;
        RECT 75.965 136.925 76.135 137.095 ;
        RECT 76.425 136.925 76.595 137.095 ;
        RECT 76.885 136.925 77.055 137.095 ;
        RECT 77.345 136.925 77.515 137.095 ;
        RECT 77.805 136.925 77.975 137.095 ;
        RECT 78.265 136.925 78.435 137.095 ;
        RECT 78.725 136.925 78.895 137.095 ;
        RECT 79.185 136.925 79.355 137.095 ;
        RECT 79.645 136.925 79.815 137.095 ;
        RECT 80.105 136.925 80.275 137.095 ;
        RECT 80.565 136.925 80.735 137.095 ;
        RECT 81.025 136.925 81.195 137.095 ;
        RECT 81.485 136.925 81.655 137.095 ;
        RECT 81.945 136.925 82.115 137.095 ;
        RECT 82.405 136.925 82.575 137.095 ;
        RECT 82.865 136.925 83.035 137.095 ;
        RECT 83.325 136.925 83.495 137.095 ;
        RECT 83.785 136.925 83.955 137.095 ;
        RECT 84.245 136.925 84.415 137.095 ;
        RECT 84.705 136.925 84.875 137.095 ;
        RECT 85.165 136.925 85.335 137.095 ;
        RECT 85.625 136.925 85.795 137.095 ;
        RECT 86.085 136.925 86.255 137.095 ;
        RECT 86.545 136.925 86.715 137.095 ;
        RECT 87.005 136.925 87.175 137.095 ;
        RECT 87.465 136.925 87.635 137.095 ;
        RECT 87.925 136.925 88.095 137.095 ;
        RECT 88.385 136.925 88.555 137.095 ;
        RECT 88.845 136.925 89.015 137.095 ;
        RECT 89.305 136.925 89.475 137.095 ;
        RECT 89.765 136.925 89.935 137.095 ;
        RECT 90.225 136.925 90.395 137.095 ;
        RECT 90.685 136.925 90.855 137.095 ;
        RECT 91.145 136.925 91.315 137.095 ;
        RECT 91.605 136.925 91.775 137.095 ;
        RECT 92.065 136.925 92.235 137.095 ;
        RECT 92.525 136.925 92.695 137.095 ;
        RECT 92.985 136.925 93.155 137.095 ;
        RECT 93.445 136.925 93.615 137.095 ;
        RECT 93.905 136.925 94.075 137.095 ;
        RECT 94.365 136.925 94.535 137.095 ;
        RECT 94.825 136.925 94.995 137.095 ;
        RECT 95.285 136.925 95.455 137.095 ;
        RECT 95.745 136.925 95.915 137.095 ;
        RECT 96.205 136.925 96.375 137.095 ;
        RECT 96.665 136.925 96.835 137.095 ;
        RECT 97.125 136.925 97.295 137.095 ;
        RECT 97.585 136.925 97.755 137.095 ;
        RECT 98.045 136.925 98.215 137.095 ;
        RECT 98.505 136.925 98.675 137.095 ;
        RECT 98.965 136.925 99.135 137.095 ;
        RECT 99.425 136.925 99.595 137.095 ;
        RECT 99.885 136.925 100.055 137.095 ;
        RECT 100.345 136.925 100.515 137.095 ;
        RECT 100.805 136.925 100.975 137.095 ;
        RECT 101.265 136.925 101.435 137.095 ;
        RECT 101.725 136.925 101.895 137.095 ;
        RECT 102.185 136.925 102.355 137.095 ;
        RECT 102.645 136.925 102.815 137.095 ;
        RECT 103.105 136.925 103.275 137.095 ;
        RECT 103.565 136.925 103.735 137.095 ;
        RECT 104.025 136.925 104.195 137.095 ;
        RECT 104.485 136.925 104.655 137.095 ;
        RECT 104.945 136.925 105.115 137.095 ;
        RECT 105.405 136.925 105.575 137.095 ;
        RECT 105.865 136.925 106.035 137.095 ;
        RECT 106.325 136.925 106.495 137.095 ;
        RECT 106.785 136.925 106.955 137.095 ;
        RECT 107.245 136.925 107.415 137.095 ;
        RECT 107.705 136.925 107.875 137.095 ;
        RECT 108.165 136.925 108.335 137.095 ;
        RECT 108.625 136.925 108.795 137.095 ;
        RECT 109.085 136.925 109.255 137.095 ;
        RECT 109.545 136.925 109.715 137.095 ;
        RECT 110.005 136.925 110.175 137.095 ;
        RECT 110.465 136.925 110.635 137.095 ;
        RECT 110.925 136.925 111.095 137.095 ;
        RECT 111.385 136.925 111.555 137.095 ;
        RECT 111.845 136.925 112.015 137.095 ;
        RECT 112.305 136.925 112.475 137.095 ;
        RECT 112.765 136.925 112.935 137.095 ;
        RECT 113.225 136.925 113.395 137.095 ;
        RECT 113.685 136.925 113.855 137.095 ;
        RECT 114.145 136.925 114.315 137.095 ;
        RECT 114.605 136.925 114.775 137.095 ;
        RECT 115.065 136.925 115.235 137.095 ;
        RECT 115.525 136.925 115.695 137.095 ;
        RECT 115.985 136.925 116.155 137.095 ;
        RECT 116.445 136.925 116.615 137.095 ;
        RECT 116.905 136.925 117.075 137.095 ;
        RECT 117.365 136.925 117.535 137.095 ;
        RECT 117.825 136.925 117.995 137.095 ;
        RECT 118.285 136.925 118.455 137.095 ;
        RECT 118.745 136.925 118.915 137.095 ;
        RECT 119.205 136.925 119.375 137.095 ;
        RECT 119.665 136.925 119.835 137.095 ;
        RECT 120.125 136.925 120.295 137.095 ;
        RECT 120.585 136.925 120.755 137.095 ;
        RECT 121.045 136.925 121.215 137.095 ;
        RECT 121.505 136.925 121.675 137.095 ;
        RECT 121.965 136.925 122.135 137.095 ;
        RECT 122.425 136.925 122.595 137.095 ;
        RECT 122.885 136.925 123.055 137.095 ;
        RECT 123.345 136.925 123.515 137.095 ;
        RECT 123.805 136.925 123.975 137.095 ;
        RECT 124.265 136.925 124.435 137.095 ;
        RECT 124.725 136.925 124.895 137.095 ;
        RECT 125.185 136.925 125.355 137.095 ;
        RECT 125.645 136.925 125.815 137.095 ;
        RECT 126.105 136.925 126.275 137.095 ;
        RECT 126.565 136.925 126.735 137.095 ;
        RECT 127.025 136.925 127.195 137.095 ;
        RECT 127.485 136.925 127.655 137.095 ;
        RECT 127.945 136.925 128.115 137.095 ;
        RECT 128.405 136.925 128.575 137.095 ;
        RECT 128.865 136.925 129.035 137.095 ;
        RECT 129.325 136.925 129.495 137.095 ;
        RECT 129.785 136.925 129.955 137.095 ;
        RECT 130.245 136.925 130.415 137.095 ;
        RECT 130.705 136.925 130.875 137.095 ;
        RECT 131.165 136.925 131.335 137.095 ;
        RECT 131.625 136.925 131.795 137.095 ;
        RECT 132.085 136.925 132.255 137.095 ;
        RECT 132.545 136.925 132.715 137.095 ;
        RECT 133.005 136.925 133.175 137.095 ;
        RECT 133.465 136.925 133.635 137.095 ;
        RECT 133.925 136.925 134.095 137.095 ;
        RECT 134.385 136.925 134.555 137.095 ;
        RECT 134.845 136.925 135.015 137.095 ;
        RECT 135.305 136.925 135.475 137.095 ;
        RECT 135.765 136.925 135.935 137.095 ;
        RECT 136.225 136.925 136.395 137.095 ;
        RECT 136.685 136.925 136.855 137.095 ;
        RECT 137.145 136.925 137.315 137.095 ;
        RECT 137.605 136.925 137.775 137.095 ;
        RECT 138.065 136.925 138.235 137.095 ;
        RECT 138.525 136.925 138.695 137.095 ;
        RECT 138.985 136.925 139.155 137.095 ;
        RECT 50.665 134.205 50.835 134.375 ;
        RECT 51.125 134.205 51.295 134.375 ;
        RECT 51.585 134.205 51.755 134.375 ;
        RECT 52.045 134.205 52.215 134.375 ;
        RECT 52.505 134.205 52.675 134.375 ;
        RECT 52.965 134.205 53.135 134.375 ;
        RECT 53.425 134.205 53.595 134.375 ;
        RECT 53.885 134.205 54.055 134.375 ;
        RECT 54.345 134.205 54.515 134.375 ;
        RECT 54.805 134.205 54.975 134.375 ;
        RECT 55.265 134.205 55.435 134.375 ;
        RECT 55.725 134.205 55.895 134.375 ;
        RECT 56.185 134.205 56.355 134.375 ;
        RECT 56.645 134.205 56.815 134.375 ;
        RECT 57.105 134.205 57.275 134.375 ;
        RECT 57.565 134.205 57.735 134.375 ;
        RECT 58.025 134.205 58.195 134.375 ;
        RECT 58.485 134.205 58.655 134.375 ;
        RECT 58.945 134.205 59.115 134.375 ;
        RECT 59.405 134.205 59.575 134.375 ;
        RECT 59.865 134.205 60.035 134.375 ;
        RECT 60.325 134.205 60.495 134.375 ;
        RECT 60.785 134.205 60.955 134.375 ;
        RECT 61.245 134.205 61.415 134.375 ;
        RECT 61.705 134.205 61.875 134.375 ;
        RECT 62.165 134.205 62.335 134.375 ;
        RECT 62.625 134.205 62.795 134.375 ;
        RECT 63.085 134.205 63.255 134.375 ;
        RECT 63.545 134.205 63.715 134.375 ;
        RECT 64.005 134.205 64.175 134.375 ;
        RECT 64.465 134.205 64.635 134.375 ;
        RECT 64.925 134.205 65.095 134.375 ;
        RECT 65.385 134.205 65.555 134.375 ;
        RECT 65.845 134.205 66.015 134.375 ;
        RECT 66.305 134.205 66.475 134.375 ;
        RECT 66.765 134.205 66.935 134.375 ;
        RECT 67.225 134.205 67.395 134.375 ;
        RECT 67.685 134.205 67.855 134.375 ;
        RECT 68.145 134.205 68.315 134.375 ;
        RECT 68.605 134.205 68.775 134.375 ;
        RECT 69.065 134.205 69.235 134.375 ;
        RECT 69.525 134.205 69.695 134.375 ;
        RECT 69.985 134.205 70.155 134.375 ;
        RECT 70.445 134.205 70.615 134.375 ;
        RECT 70.905 134.205 71.075 134.375 ;
        RECT 71.365 134.205 71.535 134.375 ;
        RECT 71.825 134.205 71.995 134.375 ;
        RECT 72.285 134.205 72.455 134.375 ;
        RECT 72.745 134.205 72.915 134.375 ;
        RECT 73.205 134.205 73.375 134.375 ;
        RECT 73.665 134.205 73.835 134.375 ;
        RECT 74.125 134.205 74.295 134.375 ;
        RECT 74.585 134.205 74.755 134.375 ;
        RECT 75.045 134.205 75.215 134.375 ;
        RECT 75.505 134.205 75.675 134.375 ;
        RECT 75.965 134.205 76.135 134.375 ;
        RECT 76.425 134.205 76.595 134.375 ;
        RECT 76.885 134.205 77.055 134.375 ;
        RECT 77.345 134.205 77.515 134.375 ;
        RECT 77.805 134.205 77.975 134.375 ;
        RECT 78.265 134.205 78.435 134.375 ;
        RECT 78.725 134.205 78.895 134.375 ;
        RECT 79.185 134.205 79.355 134.375 ;
        RECT 79.645 134.205 79.815 134.375 ;
        RECT 80.105 134.205 80.275 134.375 ;
        RECT 80.565 134.205 80.735 134.375 ;
        RECT 81.025 134.205 81.195 134.375 ;
        RECT 81.485 134.205 81.655 134.375 ;
        RECT 81.945 134.205 82.115 134.375 ;
        RECT 82.405 134.205 82.575 134.375 ;
        RECT 82.865 134.205 83.035 134.375 ;
        RECT 83.325 134.205 83.495 134.375 ;
        RECT 83.785 134.205 83.955 134.375 ;
        RECT 84.245 134.205 84.415 134.375 ;
        RECT 84.705 134.205 84.875 134.375 ;
        RECT 85.165 134.205 85.335 134.375 ;
        RECT 85.625 134.205 85.795 134.375 ;
        RECT 86.085 134.205 86.255 134.375 ;
        RECT 86.545 134.205 86.715 134.375 ;
        RECT 87.005 134.205 87.175 134.375 ;
        RECT 87.465 134.205 87.635 134.375 ;
        RECT 87.925 134.205 88.095 134.375 ;
        RECT 88.385 134.205 88.555 134.375 ;
        RECT 88.845 134.205 89.015 134.375 ;
        RECT 89.305 134.205 89.475 134.375 ;
        RECT 89.765 134.205 89.935 134.375 ;
        RECT 90.225 134.205 90.395 134.375 ;
        RECT 90.685 134.205 90.855 134.375 ;
        RECT 91.145 134.205 91.315 134.375 ;
        RECT 91.605 134.205 91.775 134.375 ;
        RECT 92.065 134.205 92.235 134.375 ;
        RECT 92.525 134.205 92.695 134.375 ;
        RECT 92.985 134.205 93.155 134.375 ;
        RECT 93.445 134.205 93.615 134.375 ;
        RECT 93.905 134.205 94.075 134.375 ;
        RECT 94.365 134.205 94.535 134.375 ;
        RECT 94.825 134.205 94.995 134.375 ;
        RECT 95.285 134.205 95.455 134.375 ;
        RECT 95.745 134.205 95.915 134.375 ;
        RECT 96.205 134.205 96.375 134.375 ;
        RECT 96.665 134.205 96.835 134.375 ;
        RECT 97.125 134.205 97.295 134.375 ;
        RECT 97.585 134.205 97.755 134.375 ;
        RECT 98.045 134.205 98.215 134.375 ;
        RECT 98.505 134.205 98.675 134.375 ;
        RECT 98.965 134.205 99.135 134.375 ;
        RECT 99.425 134.205 99.595 134.375 ;
        RECT 99.885 134.205 100.055 134.375 ;
        RECT 100.345 134.205 100.515 134.375 ;
        RECT 100.805 134.205 100.975 134.375 ;
        RECT 101.265 134.205 101.435 134.375 ;
        RECT 101.725 134.205 101.895 134.375 ;
        RECT 102.185 134.205 102.355 134.375 ;
        RECT 102.645 134.205 102.815 134.375 ;
        RECT 103.105 134.205 103.275 134.375 ;
        RECT 103.565 134.205 103.735 134.375 ;
        RECT 104.025 134.205 104.195 134.375 ;
        RECT 104.485 134.205 104.655 134.375 ;
        RECT 104.945 134.205 105.115 134.375 ;
        RECT 105.405 134.205 105.575 134.375 ;
        RECT 105.865 134.205 106.035 134.375 ;
        RECT 106.325 134.205 106.495 134.375 ;
        RECT 106.785 134.205 106.955 134.375 ;
        RECT 107.245 134.205 107.415 134.375 ;
        RECT 107.705 134.205 107.875 134.375 ;
        RECT 108.165 134.205 108.335 134.375 ;
        RECT 108.625 134.205 108.795 134.375 ;
        RECT 109.085 134.205 109.255 134.375 ;
        RECT 109.545 134.205 109.715 134.375 ;
        RECT 110.005 134.205 110.175 134.375 ;
        RECT 110.465 134.205 110.635 134.375 ;
        RECT 110.925 134.205 111.095 134.375 ;
        RECT 111.385 134.205 111.555 134.375 ;
        RECT 111.845 134.205 112.015 134.375 ;
        RECT 112.305 134.205 112.475 134.375 ;
        RECT 112.765 134.205 112.935 134.375 ;
        RECT 113.225 134.205 113.395 134.375 ;
        RECT 113.685 134.205 113.855 134.375 ;
        RECT 114.145 134.205 114.315 134.375 ;
        RECT 114.605 134.205 114.775 134.375 ;
        RECT 115.065 134.205 115.235 134.375 ;
        RECT 115.525 134.205 115.695 134.375 ;
        RECT 115.985 134.205 116.155 134.375 ;
        RECT 116.445 134.205 116.615 134.375 ;
        RECT 116.905 134.205 117.075 134.375 ;
        RECT 117.365 134.205 117.535 134.375 ;
        RECT 117.825 134.205 117.995 134.375 ;
        RECT 118.285 134.205 118.455 134.375 ;
        RECT 118.745 134.205 118.915 134.375 ;
        RECT 119.205 134.205 119.375 134.375 ;
        RECT 119.665 134.205 119.835 134.375 ;
        RECT 120.125 134.205 120.295 134.375 ;
        RECT 120.585 134.205 120.755 134.375 ;
        RECT 121.045 134.205 121.215 134.375 ;
        RECT 121.505 134.205 121.675 134.375 ;
        RECT 121.965 134.205 122.135 134.375 ;
        RECT 122.425 134.205 122.595 134.375 ;
        RECT 122.885 134.205 123.055 134.375 ;
        RECT 123.345 134.205 123.515 134.375 ;
        RECT 123.805 134.205 123.975 134.375 ;
        RECT 124.265 134.205 124.435 134.375 ;
        RECT 124.725 134.205 124.895 134.375 ;
        RECT 125.185 134.205 125.355 134.375 ;
        RECT 125.645 134.205 125.815 134.375 ;
        RECT 126.105 134.205 126.275 134.375 ;
        RECT 126.565 134.205 126.735 134.375 ;
        RECT 127.025 134.205 127.195 134.375 ;
        RECT 127.485 134.205 127.655 134.375 ;
        RECT 127.945 134.205 128.115 134.375 ;
        RECT 128.405 134.205 128.575 134.375 ;
        RECT 128.865 134.205 129.035 134.375 ;
        RECT 129.325 134.205 129.495 134.375 ;
        RECT 129.785 134.205 129.955 134.375 ;
        RECT 130.245 134.205 130.415 134.375 ;
        RECT 130.705 134.205 130.875 134.375 ;
        RECT 131.165 134.205 131.335 134.375 ;
        RECT 131.625 134.205 131.795 134.375 ;
        RECT 132.085 134.205 132.255 134.375 ;
        RECT 132.545 134.205 132.715 134.375 ;
        RECT 133.005 134.205 133.175 134.375 ;
        RECT 133.465 134.205 133.635 134.375 ;
        RECT 133.925 134.205 134.095 134.375 ;
        RECT 134.385 134.205 134.555 134.375 ;
        RECT 134.845 134.205 135.015 134.375 ;
        RECT 135.305 134.205 135.475 134.375 ;
        RECT 135.765 134.205 135.935 134.375 ;
        RECT 136.225 134.205 136.395 134.375 ;
        RECT 136.685 134.205 136.855 134.375 ;
        RECT 137.145 134.205 137.315 134.375 ;
        RECT 137.605 134.205 137.775 134.375 ;
        RECT 138.065 134.205 138.235 134.375 ;
        RECT 138.525 134.205 138.695 134.375 ;
        RECT 138.985 134.205 139.155 134.375 ;
        RECT 50.665 131.485 50.835 131.655 ;
        RECT 51.125 131.485 51.295 131.655 ;
        RECT 51.585 131.485 51.755 131.655 ;
        RECT 52.045 131.485 52.215 131.655 ;
        RECT 52.505 131.485 52.675 131.655 ;
        RECT 52.965 131.485 53.135 131.655 ;
        RECT 53.425 131.485 53.595 131.655 ;
        RECT 53.885 131.485 54.055 131.655 ;
        RECT 54.345 131.485 54.515 131.655 ;
        RECT 54.805 131.485 54.975 131.655 ;
        RECT 55.265 131.485 55.435 131.655 ;
        RECT 55.725 131.485 55.895 131.655 ;
        RECT 56.185 131.485 56.355 131.655 ;
        RECT 56.645 131.485 56.815 131.655 ;
        RECT 57.105 131.485 57.275 131.655 ;
        RECT 57.565 131.485 57.735 131.655 ;
        RECT 58.025 131.485 58.195 131.655 ;
        RECT 58.485 131.485 58.655 131.655 ;
        RECT 58.945 131.485 59.115 131.655 ;
        RECT 59.405 131.485 59.575 131.655 ;
        RECT 59.865 131.485 60.035 131.655 ;
        RECT 60.325 131.485 60.495 131.655 ;
        RECT 60.785 131.485 60.955 131.655 ;
        RECT 61.245 131.485 61.415 131.655 ;
        RECT 61.705 131.485 61.875 131.655 ;
        RECT 62.165 131.485 62.335 131.655 ;
        RECT 62.625 131.485 62.795 131.655 ;
        RECT 63.085 131.485 63.255 131.655 ;
        RECT 63.545 131.485 63.715 131.655 ;
        RECT 64.005 131.485 64.175 131.655 ;
        RECT 64.465 131.485 64.635 131.655 ;
        RECT 64.925 131.485 65.095 131.655 ;
        RECT 65.385 131.485 65.555 131.655 ;
        RECT 65.845 131.485 66.015 131.655 ;
        RECT 66.305 131.485 66.475 131.655 ;
        RECT 66.765 131.485 66.935 131.655 ;
        RECT 67.225 131.485 67.395 131.655 ;
        RECT 67.685 131.485 67.855 131.655 ;
        RECT 68.145 131.485 68.315 131.655 ;
        RECT 68.605 131.485 68.775 131.655 ;
        RECT 69.065 131.485 69.235 131.655 ;
        RECT 69.525 131.485 69.695 131.655 ;
        RECT 69.985 131.485 70.155 131.655 ;
        RECT 70.445 131.485 70.615 131.655 ;
        RECT 70.905 131.485 71.075 131.655 ;
        RECT 71.365 131.485 71.535 131.655 ;
        RECT 71.825 131.485 71.995 131.655 ;
        RECT 72.285 131.485 72.455 131.655 ;
        RECT 72.745 131.485 72.915 131.655 ;
        RECT 73.205 131.485 73.375 131.655 ;
        RECT 73.665 131.485 73.835 131.655 ;
        RECT 74.125 131.485 74.295 131.655 ;
        RECT 74.585 131.485 74.755 131.655 ;
        RECT 75.045 131.485 75.215 131.655 ;
        RECT 75.505 131.485 75.675 131.655 ;
        RECT 75.965 131.485 76.135 131.655 ;
        RECT 76.425 131.485 76.595 131.655 ;
        RECT 76.885 131.485 77.055 131.655 ;
        RECT 77.345 131.485 77.515 131.655 ;
        RECT 77.805 131.485 77.975 131.655 ;
        RECT 78.265 131.485 78.435 131.655 ;
        RECT 78.725 131.485 78.895 131.655 ;
        RECT 79.185 131.485 79.355 131.655 ;
        RECT 79.645 131.485 79.815 131.655 ;
        RECT 80.105 131.485 80.275 131.655 ;
        RECT 80.565 131.485 80.735 131.655 ;
        RECT 81.025 131.485 81.195 131.655 ;
        RECT 81.485 131.485 81.655 131.655 ;
        RECT 81.945 131.485 82.115 131.655 ;
        RECT 82.405 131.485 82.575 131.655 ;
        RECT 82.865 131.485 83.035 131.655 ;
        RECT 83.325 131.485 83.495 131.655 ;
        RECT 83.785 131.485 83.955 131.655 ;
        RECT 84.245 131.485 84.415 131.655 ;
        RECT 84.705 131.485 84.875 131.655 ;
        RECT 85.165 131.485 85.335 131.655 ;
        RECT 85.625 131.485 85.795 131.655 ;
        RECT 86.085 131.485 86.255 131.655 ;
        RECT 86.545 131.485 86.715 131.655 ;
        RECT 87.005 131.485 87.175 131.655 ;
        RECT 87.465 131.485 87.635 131.655 ;
        RECT 87.925 131.485 88.095 131.655 ;
        RECT 88.385 131.485 88.555 131.655 ;
        RECT 88.845 131.485 89.015 131.655 ;
        RECT 89.305 131.485 89.475 131.655 ;
        RECT 89.765 131.485 89.935 131.655 ;
        RECT 90.225 131.485 90.395 131.655 ;
        RECT 90.685 131.485 90.855 131.655 ;
        RECT 91.145 131.485 91.315 131.655 ;
        RECT 91.605 131.485 91.775 131.655 ;
        RECT 92.065 131.485 92.235 131.655 ;
        RECT 92.525 131.485 92.695 131.655 ;
        RECT 92.985 131.485 93.155 131.655 ;
        RECT 93.445 131.485 93.615 131.655 ;
        RECT 93.905 131.485 94.075 131.655 ;
        RECT 94.365 131.485 94.535 131.655 ;
        RECT 94.825 131.485 94.995 131.655 ;
        RECT 95.285 131.485 95.455 131.655 ;
        RECT 95.745 131.485 95.915 131.655 ;
        RECT 96.205 131.485 96.375 131.655 ;
        RECT 96.665 131.485 96.835 131.655 ;
        RECT 97.125 131.485 97.295 131.655 ;
        RECT 97.585 131.485 97.755 131.655 ;
        RECT 98.045 131.485 98.215 131.655 ;
        RECT 98.505 131.485 98.675 131.655 ;
        RECT 98.965 131.485 99.135 131.655 ;
        RECT 99.425 131.485 99.595 131.655 ;
        RECT 99.885 131.485 100.055 131.655 ;
        RECT 100.345 131.485 100.515 131.655 ;
        RECT 100.805 131.485 100.975 131.655 ;
        RECT 101.265 131.485 101.435 131.655 ;
        RECT 101.725 131.485 101.895 131.655 ;
        RECT 102.185 131.485 102.355 131.655 ;
        RECT 102.645 131.485 102.815 131.655 ;
        RECT 103.105 131.485 103.275 131.655 ;
        RECT 103.565 131.485 103.735 131.655 ;
        RECT 104.025 131.485 104.195 131.655 ;
        RECT 104.485 131.485 104.655 131.655 ;
        RECT 104.945 131.485 105.115 131.655 ;
        RECT 105.405 131.485 105.575 131.655 ;
        RECT 105.865 131.485 106.035 131.655 ;
        RECT 106.325 131.485 106.495 131.655 ;
        RECT 106.785 131.485 106.955 131.655 ;
        RECT 107.245 131.485 107.415 131.655 ;
        RECT 107.705 131.485 107.875 131.655 ;
        RECT 108.165 131.485 108.335 131.655 ;
        RECT 108.625 131.485 108.795 131.655 ;
        RECT 109.085 131.485 109.255 131.655 ;
        RECT 109.545 131.485 109.715 131.655 ;
        RECT 110.005 131.485 110.175 131.655 ;
        RECT 110.465 131.485 110.635 131.655 ;
        RECT 110.925 131.485 111.095 131.655 ;
        RECT 111.385 131.485 111.555 131.655 ;
        RECT 111.845 131.485 112.015 131.655 ;
        RECT 112.305 131.485 112.475 131.655 ;
        RECT 112.765 131.485 112.935 131.655 ;
        RECT 113.225 131.485 113.395 131.655 ;
        RECT 113.685 131.485 113.855 131.655 ;
        RECT 114.145 131.485 114.315 131.655 ;
        RECT 114.605 131.485 114.775 131.655 ;
        RECT 115.065 131.485 115.235 131.655 ;
        RECT 115.525 131.485 115.695 131.655 ;
        RECT 115.985 131.485 116.155 131.655 ;
        RECT 116.445 131.485 116.615 131.655 ;
        RECT 116.905 131.485 117.075 131.655 ;
        RECT 117.365 131.485 117.535 131.655 ;
        RECT 117.825 131.485 117.995 131.655 ;
        RECT 118.285 131.485 118.455 131.655 ;
        RECT 118.745 131.485 118.915 131.655 ;
        RECT 119.205 131.485 119.375 131.655 ;
        RECT 119.665 131.485 119.835 131.655 ;
        RECT 120.125 131.485 120.295 131.655 ;
        RECT 120.585 131.485 120.755 131.655 ;
        RECT 121.045 131.485 121.215 131.655 ;
        RECT 121.505 131.485 121.675 131.655 ;
        RECT 121.965 131.485 122.135 131.655 ;
        RECT 122.425 131.485 122.595 131.655 ;
        RECT 122.885 131.485 123.055 131.655 ;
        RECT 123.345 131.485 123.515 131.655 ;
        RECT 123.805 131.485 123.975 131.655 ;
        RECT 124.265 131.485 124.435 131.655 ;
        RECT 124.725 131.485 124.895 131.655 ;
        RECT 125.185 131.485 125.355 131.655 ;
        RECT 125.645 131.485 125.815 131.655 ;
        RECT 126.105 131.485 126.275 131.655 ;
        RECT 126.565 131.485 126.735 131.655 ;
        RECT 127.025 131.485 127.195 131.655 ;
        RECT 127.485 131.485 127.655 131.655 ;
        RECT 127.945 131.485 128.115 131.655 ;
        RECT 128.405 131.485 128.575 131.655 ;
        RECT 128.865 131.485 129.035 131.655 ;
        RECT 129.325 131.485 129.495 131.655 ;
        RECT 129.785 131.485 129.955 131.655 ;
        RECT 130.245 131.485 130.415 131.655 ;
        RECT 130.705 131.485 130.875 131.655 ;
        RECT 131.165 131.485 131.335 131.655 ;
        RECT 131.625 131.485 131.795 131.655 ;
        RECT 132.085 131.485 132.255 131.655 ;
        RECT 132.545 131.485 132.715 131.655 ;
        RECT 133.005 131.485 133.175 131.655 ;
        RECT 133.465 131.485 133.635 131.655 ;
        RECT 133.925 131.485 134.095 131.655 ;
        RECT 134.385 131.485 134.555 131.655 ;
        RECT 134.845 131.485 135.015 131.655 ;
        RECT 135.305 131.485 135.475 131.655 ;
        RECT 135.765 131.485 135.935 131.655 ;
        RECT 136.225 131.485 136.395 131.655 ;
        RECT 136.685 131.485 136.855 131.655 ;
        RECT 137.145 131.485 137.315 131.655 ;
        RECT 137.605 131.485 137.775 131.655 ;
        RECT 138.065 131.485 138.235 131.655 ;
        RECT 138.525 131.485 138.695 131.655 ;
        RECT 138.985 131.485 139.155 131.655 ;
        RECT 50.665 128.765 50.835 128.935 ;
        RECT 51.125 128.765 51.295 128.935 ;
        RECT 51.585 128.765 51.755 128.935 ;
        RECT 52.045 128.765 52.215 128.935 ;
        RECT 52.505 128.765 52.675 128.935 ;
        RECT 52.965 128.765 53.135 128.935 ;
        RECT 53.425 128.765 53.595 128.935 ;
        RECT 53.885 128.765 54.055 128.935 ;
        RECT 54.345 128.765 54.515 128.935 ;
        RECT 54.805 128.765 54.975 128.935 ;
        RECT 55.265 128.765 55.435 128.935 ;
        RECT 55.725 128.765 55.895 128.935 ;
        RECT 56.185 128.765 56.355 128.935 ;
        RECT 56.645 128.765 56.815 128.935 ;
        RECT 57.105 128.765 57.275 128.935 ;
        RECT 57.565 128.765 57.735 128.935 ;
        RECT 58.025 128.765 58.195 128.935 ;
        RECT 58.485 128.765 58.655 128.935 ;
        RECT 58.945 128.765 59.115 128.935 ;
        RECT 59.405 128.765 59.575 128.935 ;
        RECT 59.865 128.765 60.035 128.935 ;
        RECT 60.325 128.765 60.495 128.935 ;
        RECT 60.785 128.765 60.955 128.935 ;
        RECT 61.245 128.765 61.415 128.935 ;
        RECT 61.705 128.765 61.875 128.935 ;
        RECT 62.165 128.765 62.335 128.935 ;
        RECT 62.625 128.765 62.795 128.935 ;
        RECT 63.085 128.765 63.255 128.935 ;
        RECT 63.545 128.765 63.715 128.935 ;
        RECT 64.005 128.765 64.175 128.935 ;
        RECT 64.465 128.765 64.635 128.935 ;
        RECT 64.925 128.765 65.095 128.935 ;
        RECT 65.385 128.765 65.555 128.935 ;
        RECT 65.845 128.765 66.015 128.935 ;
        RECT 66.305 128.765 66.475 128.935 ;
        RECT 66.765 128.765 66.935 128.935 ;
        RECT 67.225 128.765 67.395 128.935 ;
        RECT 67.685 128.765 67.855 128.935 ;
        RECT 68.145 128.765 68.315 128.935 ;
        RECT 68.605 128.765 68.775 128.935 ;
        RECT 69.065 128.765 69.235 128.935 ;
        RECT 69.525 128.765 69.695 128.935 ;
        RECT 69.985 128.765 70.155 128.935 ;
        RECT 70.445 128.765 70.615 128.935 ;
        RECT 70.905 128.765 71.075 128.935 ;
        RECT 71.365 128.765 71.535 128.935 ;
        RECT 71.825 128.765 71.995 128.935 ;
        RECT 72.285 128.765 72.455 128.935 ;
        RECT 72.745 128.765 72.915 128.935 ;
        RECT 73.205 128.765 73.375 128.935 ;
        RECT 73.665 128.765 73.835 128.935 ;
        RECT 74.125 128.765 74.295 128.935 ;
        RECT 74.585 128.765 74.755 128.935 ;
        RECT 75.045 128.765 75.215 128.935 ;
        RECT 75.505 128.765 75.675 128.935 ;
        RECT 75.965 128.765 76.135 128.935 ;
        RECT 76.425 128.765 76.595 128.935 ;
        RECT 76.885 128.765 77.055 128.935 ;
        RECT 77.345 128.765 77.515 128.935 ;
        RECT 77.805 128.765 77.975 128.935 ;
        RECT 78.265 128.765 78.435 128.935 ;
        RECT 78.725 128.765 78.895 128.935 ;
        RECT 79.185 128.765 79.355 128.935 ;
        RECT 79.645 128.765 79.815 128.935 ;
        RECT 80.105 128.765 80.275 128.935 ;
        RECT 80.565 128.765 80.735 128.935 ;
        RECT 81.025 128.765 81.195 128.935 ;
        RECT 81.485 128.765 81.655 128.935 ;
        RECT 81.945 128.765 82.115 128.935 ;
        RECT 82.405 128.765 82.575 128.935 ;
        RECT 82.865 128.765 83.035 128.935 ;
        RECT 83.325 128.765 83.495 128.935 ;
        RECT 83.785 128.765 83.955 128.935 ;
        RECT 84.245 128.765 84.415 128.935 ;
        RECT 84.705 128.765 84.875 128.935 ;
        RECT 85.165 128.765 85.335 128.935 ;
        RECT 85.625 128.765 85.795 128.935 ;
        RECT 86.085 128.765 86.255 128.935 ;
        RECT 86.545 128.765 86.715 128.935 ;
        RECT 87.005 128.765 87.175 128.935 ;
        RECT 87.465 128.765 87.635 128.935 ;
        RECT 87.925 128.765 88.095 128.935 ;
        RECT 88.385 128.765 88.555 128.935 ;
        RECT 88.845 128.765 89.015 128.935 ;
        RECT 89.305 128.765 89.475 128.935 ;
        RECT 89.765 128.765 89.935 128.935 ;
        RECT 90.225 128.765 90.395 128.935 ;
        RECT 90.685 128.765 90.855 128.935 ;
        RECT 91.145 128.765 91.315 128.935 ;
        RECT 91.605 128.765 91.775 128.935 ;
        RECT 92.065 128.765 92.235 128.935 ;
        RECT 92.525 128.765 92.695 128.935 ;
        RECT 92.985 128.765 93.155 128.935 ;
        RECT 93.445 128.765 93.615 128.935 ;
        RECT 93.905 128.765 94.075 128.935 ;
        RECT 94.365 128.765 94.535 128.935 ;
        RECT 94.825 128.765 94.995 128.935 ;
        RECT 95.285 128.765 95.455 128.935 ;
        RECT 95.745 128.765 95.915 128.935 ;
        RECT 96.205 128.765 96.375 128.935 ;
        RECT 96.665 128.765 96.835 128.935 ;
        RECT 97.125 128.765 97.295 128.935 ;
        RECT 97.585 128.765 97.755 128.935 ;
        RECT 98.045 128.765 98.215 128.935 ;
        RECT 98.505 128.765 98.675 128.935 ;
        RECT 98.965 128.765 99.135 128.935 ;
        RECT 99.425 128.765 99.595 128.935 ;
        RECT 99.885 128.765 100.055 128.935 ;
        RECT 100.345 128.765 100.515 128.935 ;
        RECT 100.805 128.765 100.975 128.935 ;
        RECT 101.265 128.765 101.435 128.935 ;
        RECT 101.725 128.765 101.895 128.935 ;
        RECT 102.185 128.765 102.355 128.935 ;
        RECT 102.645 128.765 102.815 128.935 ;
        RECT 103.105 128.765 103.275 128.935 ;
        RECT 103.565 128.765 103.735 128.935 ;
        RECT 104.025 128.765 104.195 128.935 ;
        RECT 104.485 128.765 104.655 128.935 ;
        RECT 104.945 128.765 105.115 128.935 ;
        RECT 105.405 128.765 105.575 128.935 ;
        RECT 105.865 128.765 106.035 128.935 ;
        RECT 106.325 128.765 106.495 128.935 ;
        RECT 106.785 128.765 106.955 128.935 ;
        RECT 107.245 128.765 107.415 128.935 ;
        RECT 107.705 128.765 107.875 128.935 ;
        RECT 108.165 128.765 108.335 128.935 ;
        RECT 108.625 128.765 108.795 128.935 ;
        RECT 109.085 128.765 109.255 128.935 ;
        RECT 109.545 128.765 109.715 128.935 ;
        RECT 110.005 128.765 110.175 128.935 ;
        RECT 110.465 128.765 110.635 128.935 ;
        RECT 110.925 128.765 111.095 128.935 ;
        RECT 111.385 128.765 111.555 128.935 ;
        RECT 111.845 128.765 112.015 128.935 ;
        RECT 112.305 128.765 112.475 128.935 ;
        RECT 112.765 128.765 112.935 128.935 ;
        RECT 113.225 128.765 113.395 128.935 ;
        RECT 113.685 128.765 113.855 128.935 ;
        RECT 114.145 128.765 114.315 128.935 ;
        RECT 114.605 128.765 114.775 128.935 ;
        RECT 115.065 128.765 115.235 128.935 ;
        RECT 115.525 128.765 115.695 128.935 ;
        RECT 115.985 128.765 116.155 128.935 ;
        RECT 116.445 128.765 116.615 128.935 ;
        RECT 116.905 128.765 117.075 128.935 ;
        RECT 117.365 128.765 117.535 128.935 ;
        RECT 117.825 128.765 117.995 128.935 ;
        RECT 118.285 128.765 118.455 128.935 ;
        RECT 118.745 128.765 118.915 128.935 ;
        RECT 119.205 128.765 119.375 128.935 ;
        RECT 119.665 128.765 119.835 128.935 ;
        RECT 120.125 128.765 120.295 128.935 ;
        RECT 120.585 128.765 120.755 128.935 ;
        RECT 121.045 128.765 121.215 128.935 ;
        RECT 121.505 128.765 121.675 128.935 ;
        RECT 121.965 128.765 122.135 128.935 ;
        RECT 122.425 128.765 122.595 128.935 ;
        RECT 122.885 128.765 123.055 128.935 ;
        RECT 123.345 128.765 123.515 128.935 ;
        RECT 123.805 128.765 123.975 128.935 ;
        RECT 124.265 128.765 124.435 128.935 ;
        RECT 124.725 128.765 124.895 128.935 ;
        RECT 125.185 128.765 125.355 128.935 ;
        RECT 125.645 128.765 125.815 128.935 ;
        RECT 126.105 128.765 126.275 128.935 ;
        RECT 126.565 128.765 126.735 128.935 ;
        RECT 127.025 128.765 127.195 128.935 ;
        RECT 127.485 128.765 127.655 128.935 ;
        RECT 127.945 128.765 128.115 128.935 ;
        RECT 128.405 128.765 128.575 128.935 ;
        RECT 128.865 128.765 129.035 128.935 ;
        RECT 129.325 128.765 129.495 128.935 ;
        RECT 129.785 128.765 129.955 128.935 ;
        RECT 130.245 128.765 130.415 128.935 ;
        RECT 130.705 128.765 130.875 128.935 ;
        RECT 131.165 128.765 131.335 128.935 ;
        RECT 131.625 128.765 131.795 128.935 ;
        RECT 132.085 128.765 132.255 128.935 ;
        RECT 132.545 128.765 132.715 128.935 ;
        RECT 133.005 128.765 133.175 128.935 ;
        RECT 133.465 128.765 133.635 128.935 ;
        RECT 133.925 128.765 134.095 128.935 ;
        RECT 134.385 128.765 134.555 128.935 ;
        RECT 134.845 128.765 135.015 128.935 ;
        RECT 135.305 128.765 135.475 128.935 ;
        RECT 135.765 128.765 135.935 128.935 ;
        RECT 136.225 128.765 136.395 128.935 ;
        RECT 136.685 128.765 136.855 128.935 ;
        RECT 137.145 128.765 137.315 128.935 ;
        RECT 137.605 128.765 137.775 128.935 ;
        RECT 138.065 128.765 138.235 128.935 ;
        RECT 138.525 128.765 138.695 128.935 ;
        RECT 138.985 128.765 139.155 128.935 ;
        RECT 50.665 126.045 50.835 126.215 ;
        RECT 51.125 126.045 51.295 126.215 ;
        RECT 51.585 126.045 51.755 126.215 ;
        RECT 52.045 126.045 52.215 126.215 ;
        RECT 52.505 126.045 52.675 126.215 ;
        RECT 52.965 126.045 53.135 126.215 ;
        RECT 53.425 126.045 53.595 126.215 ;
        RECT 53.885 126.045 54.055 126.215 ;
        RECT 54.345 126.045 54.515 126.215 ;
        RECT 54.805 126.045 54.975 126.215 ;
        RECT 55.265 126.045 55.435 126.215 ;
        RECT 55.725 126.045 55.895 126.215 ;
        RECT 56.185 126.045 56.355 126.215 ;
        RECT 56.645 126.045 56.815 126.215 ;
        RECT 57.105 126.045 57.275 126.215 ;
        RECT 57.565 126.045 57.735 126.215 ;
        RECT 58.025 126.045 58.195 126.215 ;
        RECT 58.485 126.045 58.655 126.215 ;
        RECT 58.945 126.045 59.115 126.215 ;
        RECT 59.405 126.045 59.575 126.215 ;
        RECT 59.865 126.045 60.035 126.215 ;
        RECT 60.325 126.045 60.495 126.215 ;
        RECT 60.785 126.045 60.955 126.215 ;
        RECT 61.245 126.045 61.415 126.215 ;
        RECT 61.705 126.045 61.875 126.215 ;
        RECT 62.165 126.045 62.335 126.215 ;
        RECT 62.625 126.045 62.795 126.215 ;
        RECT 63.085 126.045 63.255 126.215 ;
        RECT 63.545 126.045 63.715 126.215 ;
        RECT 64.005 126.045 64.175 126.215 ;
        RECT 64.465 126.045 64.635 126.215 ;
        RECT 64.925 126.045 65.095 126.215 ;
        RECT 65.385 126.045 65.555 126.215 ;
        RECT 65.845 126.045 66.015 126.215 ;
        RECT 66.305 126.045 66.475 126.215 ;
        RECT 66.765 126.045 66.935 126.215 ;
        RECT 67.225 126.045 67.395 126.215 ;
        RECT 67.685 126.045 67.855 126.215 ;
        RECT 68.145 126.045 68.315 126.215 ;
        RECT 68.605 126.045 68.775 126.215 ;
        RECT 69.065 126.045 69.235 126.215 ;
        RECT 69.525 126.045 69.695 126.215 ;
        RECT 69.985 126.045 70.155 126.215 ;
        RECT 70.445 126.045 70.615 126.215 ;
        RECT 70.905 126.045 71.075 126.215 ;
        RECT 71.365 126.045 71.535 126.215 ;
        RECT 71.825 126.045 71.995 126.215 ;
        RECT 72.285 126.045 72.455 126.215 ;
        RECT 72.745 126.045 72.915 126.215 ;
        RECT 73.205 126.045 73.375 126.215 ;
        RECT 73.665 126.045 73.835 126.215 ;
        RECT 74.125 126.045 74.295 126.215 ;
        RECT 74.585 126.045 74.755 126.215 ;
        RECT 75.045 126.045 75.215 126.215 ;
        RECT 75.505 126.045 75.675 126.215 ;
        RECT 75.965 126.045 76.135 126.215 ;
        RECT 76.425 126.045 76.595 126.215 ;
        RECT 76.885 126.045 77.055 126.215 ;
        RECT 77.345 126.045 77.515 126.215 ;
        RECT 77.805 126.045 77.975 126.215 ;
        RECT 78.265 126.045 78.435 126.215 ;
        RECT 78.725 126.045 78.895 126.215 ;
        RECT 79.185 126.045 79.355 126.215 ;
        RECT 79.645 126.045 79.815 126.215 ;
        RECT 80.105 126.045 80.275 126.215 ;
        RECT 80.565 126.045 80.735 126.215 ;
        RECT 81.025 126.045 81.195 126.215 ;
        RECT 81.485 126.045 81.655 126.215 ;
        RECT 81.945 126.045 82.115 126.215 ;
        RECT 82.405 126.045 82.575 126.215 ;
        RECT 82.865 126.045 83.035 126.215 ;
        RECT 83.325 126.045 83.495 126.215 ;
        RECT 83.785 126.045 83.955 126.215 ;
        RECT 84.245 126.045 84.415 126.215 ;
        RECT 84.705 126.045 84.875 126.215 ;
        RECT 85.165 126.045 85.335 126.215 ;
        RECT 85.625 126.045 85.795 126.215 ;
        RECT 86.085 126.045 86.255 126.215 ;
        RECT 86.545 126.045 86.715 126.215 ;
        RECT 87.005 126.045 87.175 126.215 ;
        RECT 87.465 126.045 87.635 126.215 ;
        RECT 87.925 126.045 88.095 126.215 ;
        RECT 88.385 126.045 88.555 126.215 ;
        RECT 88.845 126.045 89.015 126.215 ;
        RECT 89.305 126.045 89.475 126.215 ;
        RECT 89.765 126.045 89.935 126.215 ;
        RECT 90.225 126.045 90.395 126.215 ;
        RECT 90.685 126.045 90.855 126.215 ;
        RECT 91.145 126.045 91.315 126.215 ;
        RECT 91.605 126.045 91.775 126.215 ;
        RECT 92.065 126.045 92.235 126.215 ;
        RECT 92.525 126.045 92.695 126.215 ;
        RECT 92.985 126.045 93.155 126.215 ;
        RECT 93.445 126.045 93.615 126.215 ;
        RECT 93.905 126.045 94.075 126.215 ;
        RECT 94.365 126.045 94.535 126.215 ;
        RECT 94.825 126.045 94.995 126.215 ;
        RECT 95.285 126.045 95.455 126.215 ;
        RECT 95.745 126.045 95.915 126.215 ;
        RECT 96.205 126.045 96.375 126.215 ;
        RECT 96.665 126.045 96.835 126.215 ;
        RECT 97.125 126.045 97.295 126.215 ;
        RECT 97.585 126.045 97.755 126.215 ;
        RECT 98.045 126.045 98.215 126.215 ;
        RECT 98.505 126.045 98.675 126.215 ;
        RECT 98.965 126.045 99.135 126.215 ;
        RECT 99.425 126.045 99.595 126.215 ;
        RECT 99.885 126.045 100.055 126.215 ;
        RECT 100.345 126.045 100.515 126.215 ;
        RECT 100.805 126.045 100.975 126.215 ;
        RECT 101.265 126.045 101.435 126.215 ;
        RECT 101.725 126.045 101.895 126.215 ;
        RECT 102.185 126.045 102.355 126.215 ;
        RECT 102.645 126.045 102.815 126.215 ;
        RECT 103.105 126.045 103.275 126.215 ;
        RECT 103.565 126.045 103.735 126.215 ;
        RECT 104.025 126.045 104.195 126.215 ;
        RECT 104.485 126.045 104.655 126.215 ;
        RECT 104.945 126.045 105.115 126.215 ;
        RECT 105.405 126.045 105.575 126.215 ;
        RECT 105.865 126.045 106.035 126.215 ;
        RECT 106.325 126.045 106.495 126.215 ;
        RECT 106.785 126.045 106.955 126.215 ;
        RECT 107.245 126.045 107.415 126.215 ;
        RECT 107.705 126.045 107.875 126.215 ;
        RECT 108.165 126.045 108.335 126.215 ;
        RECT 108.625 126.045 108.795 126.215 ;
        RECT 109.085 126.045 109.255 126.215 ;
        RECT 109.545 126.045 109.715 126.215 ;
        RECT 110.005 126.045 110.175 126.215 ;
        RECT 110.465 126.045 110.635 126.215 ;
        RECT 110.925 126.045 111.095 126.215 ;
        RECT 111.385 126.045 111.555 126.215 ;
        RECT 111.845 126.045 112.015 126.215 ;
        RECT 112.305 126.045 112.475 126.215 ;
        RECT 112.765 126.045 112.935 126.215 ;
        RECT 113.225 126.045 113.395 126.215 ;
        RECT 113.685 126.045 113.855 126.215 ;
        RECT 114.145 126.045 114.315 126.215 ;
        RECT 114.605 126.045 114.775 126.215 ;
        RECT 115.065 126.045 115.235 126.215 ;
        RECT 115.525 126.045 115.695 126.215 ;
        RECT 115.985 126.045 116.155 126.215 ;
        RECT 116.445 126.045 116.615 126.215 ;
        RECT 116.905 126.045 117.075 126.215 ;
        RECT 117.365 126.045 117.535 126.215 ;
        RECT 117.825 126.045 117.995 126.215 ;
        RECT 118.285 126.045 118.455 126.215 ;
        RECT 118.745 126.045 118.915 126.215 ;
        RECT 119.205 126.045 119.375 126.215 ;
        RECT 119.665 126.045 119.835 126.215 ;
        RECT 120.125 126.045 120.295 126.215 ;
        RECT 120.585 126.045 120.755 126.215 ;
        RECT 121.045 126.045 121.215 126.215 ;
        RECT 121.505 126.045 121.675 126.215 ;
        RECT 121.965 126.045 122.135 126.215 ;
        RECT 122.425 126.045 122.595 126.215 ;
        RECT 122.885 126.045 123.055 126.215 ;
        RECT 123.345 126.045 123.515 126.215 ;
        RECT 123.805 126.045 123.975 126.215 ;
        RECT 124.265 126.045 124.435 126.215 ;
        RECT 124.725 126.045 124.895 126.215 ;
        RECT 125.185 126.045 125.355 126.215 ;
        RECT 125.645 126.045 125.815 126.215 ;
        RECT 126.105 126.045 126.275 126.215 ;
        RECT 126.565 126.045 126.735 126.215 ;
        RECT 127.025 126.045 127.195 126.215 ;
        RECT 127.485 126.045 127.655 126.215 ;
        RECT 127.945 126.045 128.115 126.215 ;
        RECT 128.405 126.045 128.575 126.215 ;
        RECT 128.865 126.045 129.035 126.215 ;
        RECT 129.325 126.045 129.495 126.215 ;
        RECT 129.785 126.045 129.955 126.215 ;
        RECT 130.245 126.045 130.415 126.215 ;
        RECT 130.705 126.045 130.875 126.215 ;
        RECT 131.165 126.045 131.335 126.215 ;
        RECT 131.625 126.045 131.795 126.215 ;
        RECT 132.085 126.045 132.255 126.215 ;
        RECT 132.545 126.045 132.715 126.215 ;
        RECT 133.005 126.045 133.175 126.215 ;
        RECT 133.465 126.045 133.635 126.215 ;
        RECT 133.925 126.045 134.095 126.215 ;
        RECT 134.385 126.045 134.555 126.215 ;
        RECT 134.845 126.045 135.015 126.215 ;
        RECT 135.305 126.045 135.475 126.215 ;
        RECT 135.765 126.045 135.935 126.215 ;
        RECT 136.225 126.045 136.395 126.215 ;
        RECT 136.685 126.045 136.855 126.215 ;
        RECT 137.145 126.045 137.315 126.215 ;
        RECT 137.605 126.045 137.775 126.215 ;
        RECT 138.065 126.045 138.235 126.215 ;
        RECT 138.525 126.045 138.695 126.215 ;
        RECT 138.985 126.045 139.155 126.215 ;
        RECT 50.665 123.325 50.835 123.495 ;
        RECT 51.125 123.325 51.295 123.495 ;
        RECT 51.585 123.325 51.755 123.495 ;
        RECT 52.045 123.325 52.215 123.495 ;
        RECT 52.505 123.325 52.675 123.495 ;
        RECT 52.965 123.325 53.135 123.495 ;
        RECT 53.425 123.325 53.595 123.495 ;
        RECT 53.885 123.325 54.055 123.495 ;
        RECT 54.345 123.325 54.515 123.495 ;
        RECT 54.805 123.325 54.975 123.495 ;
        RECT 55.265 123.325 55.435 123.495 ;
        RECT 55.725 123.325 55.895 123.495 ;
        RECT 56.185 123.325 56.355 123.495 ;
        RECT 56.645 123.325 56.815 123.495 ;
        RECT 57.105 123.325 57.275 123.495 ;
        RECT 57.565 123.325 57.735 123.495 ;
        RECT 58.025 123.325 58.195 123.495 ;
        RECT 58.485 123.325 58.655 123.495 ;
        RECT 58.945 123.325 59.115 123.495 ;
        RECT 59.405 123.325 59.575 123.495 ;
        RECT 59.865 123.325 60.035 123.495 ;
        RECT 60.325 123.325 60.495 123.495 ;
        RECT 60.785 123.325 60.955 123.495 ;
        RECT 61.245 123.325 61.415 123.495 ;
        RECT 61.705 123.325 61.875 123.495 ;
        RECT 62.165 123.325 62.335 123.495 ;
        RECT 62.625 123.325 62.795 123.495 ;
        RECT 63.085 123.325 63.255 123.495 ;
        RECT 63.545 123.325 63.715 123.495 ;
        RECT 64.005 123.325 64.175 123.495 ;
        RECT 64.465 123.325 64.635 123.495 ;
        RECT 64.925 123.325 65.095 123.495 ;
        RECT 65.385 123.325 65.555 123.495 ;
        RECT 65.845 123.325 66.015 123.495 ;
        RECT 66.305 123.325 66.475 123.495 ;
        RECT 66.765 123.325 66.935 123.495 ;
        RECT 67.225 123.325 67.395 123.495 ;
        RECT 67.685 123.325 67.855 123.495 ;
        RECT 68.145 123.325 68.315 123.495 ;
        RECT 68.605 123.325 68.775 123.495 ;
        RECT 69.065 123.325 69.235 123.495 ;
        RECT 69.525 123.325 69.695 123.495 ;
        RECT 69.985 123.325 70.155 123.495 ;
        RECT 70.445 123.325 70.615 123.495 ;
        RECT 70.905 123.325 71.075 123.495 ;
        RECT 71.365 123.325 71.535 123.495 ;
        RECT 71.825 123.325 71.995 123.495 ;
        RECT 72.285 123.325 72.455 123.495 ;
        RECT 72.745 123.325 72.915 123.495 ;
        RECT 73.205 123.325 73.375 123.495 ;
        RECT 73.665 123.325 73.835 123.495 ;
        RECT 74.125 123.325 74.295 123.495 ;
        RECT 74.585 123.325 74.755 123.495 ;
        RECT 75.045 123.325 75.215 123.495 ;
        RECT 75.505 123.325 75.675 123.495 ;
        RECT 75.965 123.325 76.135 123.495 ;
        RECT 76.425 123.325 76.595 123.495 ;
        RECT 76.885 123.325 77.055 123.495 ;
        RECT 77.345 123.325 77.515 123.495 ;
        RECT 77.805 123.325 77.975 123.495 ;
        RECT 78.265 123.325 78.435 123.495 ;
        RECT 78.725 123.325 78.895 123.495 ;
        RECT 79.185 123.325 79.355 123.495 ;
        RECT 79.645 123.325 79.815 123.495 ;
        RECT 80.105 123.325 80.275 123.495 ;
        RECT 80.565 123.325 80.735 123.495 ;
        RECT 81.025 123.325 81.195 123.495 ;
        RECT 81.485 123.325 81.655 123.495 ;
        RECT 81.945 123.325 82.115 123.495 ;
        RECT 82.405 123.325 82.575 123.495 ;
        RECT 82.865 123.325 83.035 123.495 ;
        RECT 83.325 123.325 83.495 123.495 ;
        RECT 83.785 123.325 83.955 123.495 ;
        RECT 84.245 123.325 84.415 123.495 ;
        RECT 84.705 123.325 84.875 123.495 ;
        RECT 85.165 123.325 85.335 123.495 ;
        RECT 85.625 123.325 85.795 123.495 ;
        RECT 86.085 123.325 86.255 123.495 ;
        RECT 86.545 123.325 86.715 123.495 ;
        RECT 87.005 123.325 87.175 123.495 ;
        RECT 87.465 123.325 87.635 123.495 ;
        RECT 87.925 123.325 88.095 123.495 ;
        RECT 88.385 123.325 88.555 123.495 ;
        RECT 88.845 123.325 89.015 123.495 ;
        RECT 89.305 123.325 89.475 123.495 ;
        RECT 89.765 123.325 89.935 123.495 ;
        RECT 90.225 123.325 90.395 123.495 ;
        RECT 90.685 123.325 90.855 123.495 ;
        RECT 91.145 123.325 91.315 123.495 ;
        RECT 91.605 123.325 91.775 123.495 ;
        RECT 92.065 123.325 92.235 123.495 ;
        RECT 92.525 123.325 92.695 123.495 ;
        RECT 92.985 123.325 93.155 123.495 ;
        RECT 93.445 123.325 93.615 123.495 ;
        RECT 93.905 123.325 94.075 123.495 ;
        RECT 94.365 123.325 94.535 123.495 ;
        RECT 94.825 123.325 94.995 123.495 ;
        RECT 95.285 123.325 95.455 123.495 ;
        RECT 95.745 123.325 95.915 123.495 ;
        RECT 96.205 123.325 96.375 123.495 ;
        RECT 96.665 123.325 96.835 123.495 ;
        RECT 97.125 123.325 97.295 123.495 ;
        RECT 97.585 123.325 97.755 123.495 ;
        RECT 98.045 123.325 98.215 123.495 ;
        RECT 98.505 123.325 98.675 123.495 ;
        RECT 98.965 123.325 99.135 123.495 ;
        RECT 99.425 123.325 99.595 123.495 ;
        RECT 99.885 123.325 100.055 123.495 ;
        RECT 100.345 123.325 100.515 123.495 ;
        RECT 100.805 123.325 100.975 123.495 ;
        RECT 101.265 123.325 101.435 123.495 ;
        RECT 101.725 123.325 101.895 123.495 ;
        RECT 102.185 123.325 102.355 123.495 ;
        RECT 102.645 123.325 102.815 123.495 ;
        RECT 103.105 123.325 103.275 123.495 ;
        RECT 103.565 123.325 103.735 123.495 ;
        RECT 104.025 123.325 104.195 123.495 ;
        RECT 104.485 123.325 104.655 123.495 ;
        RECT 104.945 123.325 105.115 123.495 ;
        RECT 105.405 123.325 105.575 123.495 ;
        RECT 105.865 123.325 106.035 123.495 ;
        RECT 106.325 123.325 106.495 123.495 ;
        RECT 106.785 123.325 106.955 123.495 ;
        RECT 107.245 123.325 107.415 123.495 ;
        RECT 107.705 123.325 107.875 123.495 ;
        RECT 108.165 123.325 108.335 123.495 ;
        RECT 108.625 123.325 108.795 123.495 ;
        RECT 109.085 123.325 109.255 123.495 ;
        RECT 109.545 123.325 109.715 123.495 ;
        RECT 110.005 123.325 110.175 123.495 ;
        RECT 110.465 123.325 110.635 123.495 ;
        RECT 110.925 123.325 111.095 123.495 ;
        RECT 111.385 123.325 111.555 123.495 ;
        RECT 111.845 123.325 112.015 123.495 ;
        RECT 112.305 123.325 112.475 123.495 ;
        RECT 112.765 123.325 112.935 123.495 ;
        RECT 113.225 123.325 113.395 123.495 ;
        RECT 113.685 123.325 113.855 123.495 ;
        RECT 114.145 123.325 114.315 123.495 ;
        RECT 114.605 123.325 114.775 123.495 ;
        RECT 115.065 123.325 115.235 123.495 ;
        RECT 115.525 123.325 115.695 123.495 ;
        RECT 115.985 123.325 116.155 123.495 ;
        RECT 116.445 123.325 116.615 123.495 ;
        RECT 116.905 123.325 117.075 123.495 ;
        RECT 117.365 123.325 117.535 123.495 ;
        RECT 117.825 123.325 117.995 123.495 ;
        RECT 118.285 123.325 118.455 123.495 ;
        RECT 118.745 123.325 118.915 123.495 ;
        RECT 119.205 123.325 119.375 123.495 ;
        RECT 119.665 123.325 119.835 123.495 ;
        RECT 120.125 123.325 120.295 123.495 ;
        RECT 120.585 123.325 120.755 123.495 ;
        RECT 121.045 123.325 121.215 123.495 ;
        RECT 121.505 123.325 121.675 123.495 ;
        RECT 121.965 123.325 122.135 123.495 ;
        RECT 122.425 123.325 122.595 123.495 ;
        RECT 122.885 123.325 123.055 123.495 ;
        RECT 123.345 123.325 123.515 123.495 ;
        RECT 123.805 123.325 123.975 123.495 ;
        RECT 124.265 123.325 124.435 123.495 ;
        RECT 124.725 123.325 124.895 123.495 ;
        RECT 125.185 123.325 125.355 123.495 ;
        RECT 125.645 123.325 125.815 123.495 ;
        RECT 126.105 123.325 126.275 123.495 ;
        RECT 126.565 123.325 126.735 123.495 ;
        RECT 127.025 123.325 127.195 123.495 ;
        RECT 127.485 123.325 127.655 123.495 ;
        RECT 127.945 123.325 128.115 123.495 ;
        RECT 128.405 123.325 128.575 123.495 ;
        RECT 128.865 123.325 129.035 123.495 ;
        RECT 129.325 123.325 129.495 123.495 ;
        RECT 129.785 123.325 129.955 123.495 ;
        RECT 130.245 123.325 130.415 123.495 ;
        RECT 130.705 123.325 130.875 123.495 ;
        RECT 131.165 123.325 131.335 123.495 ;
        RECT 131.625 123.325 131.795 123.495 ;
        RECT 132.085 123.325 132.255 123.495 ;
        RECT 132.545 123.325 132.715 123.495 ;
        RECT 133.005 123.325 133.175 123.495 ;
        RECT 133.465 123.325 133.635 123.495 ;
        RECT 133.925 123.325 134.095 123.495 ;
        RECT 134.385 123.325 134.555 123.495 ;
        RECT 134.845 123.325 135.015 123.495 ;
        RECT 135.305 123.325 135.475 123.495 ;
        RECT 135.765 123.325 135.935 123.495 ;
        RECT 136.225 123.325 136.395 123.495 ;
        RECT 136.685 123.325 136.855 123.495 ;
        RECT 137.145 123.325 137.315 123.495 ;
        RECT 137.605 123.325 137.775 123.495 ;
        RECT 138.065 123.325 138.235 123.495 ;
        RECT 138.525 123.325 138.695 123.495 ;
        RECT 138.985 123.325 139.155 123.495 ;
        RECT 50.665 120.605 50.835 120.775 ;
        RECT 51.125 120.605 51.295 120.775 ;
        RECT 51.585 120.605 51.755 120.775 ;
        RECT 52.045 120.605 52.215 120.775 ;
        RECT 52.505 120.605 52.675 120.775 ;
        RECT 52.965 120.605 53.135 120.775 ;
        RECT 53.425 120.605 53.595 120.775 ;
        RECT 53.885 120.605 54.055 120.775 ;
        RECT 54.345 120.605 54.515 120.775 ;
        RECT 54.805 120.605 54.975 120.775 ;
        RECT 55.265 120.605 55.435 120.775 ;
        RECT 55.725 120.605 55.895 120.775 ;
        RECT 56.185 120.605 56.355 120.775 ;
        RECT 56.645 120.605 56.815 120.775 ;
        RECT 57.105 120.605 57.275 120.775 ;
        RECT 57.565 120.605 57.735 120.775 ;
        RECT 58.025 120.605 58.195 120.775 ;
        RECT 58.485 120.605 58.655 120.775 ;
        RECT 58.945 120.605 59.115 120.775 ;
        RECT 59.405 120.605 59.575 120.775 ;
        RECT 59.865 120.605 60.035 120.775 ;
        RECT 60.325 120.605 60.495 120.775 ;
        RECT 60.785 120.605 60.955 120.775 ;
        RECT 61.245 120.605 61.415 120.775 ;
        RECT 61.705 120.605 61.875 120.775 ;
        RECT 62.165 120.605 62.335 120.775 ;
        RECT 62.625 120.605 62.795 120.775 ;
        RECT 63.085 120.605 63.255 120.775 ;
        RECT 63.545 120.605 63.715 120.775 ;
        RECT 64.005 120.605 64.175 120.775 ;
        RECT 64.465 120.605 64.635 120.775 ;
        RECT 64.925 120.605 65.095 120.775 ;
        RECT 65.385 120.605 65.555 120.775 ;
        RECT 65.845 120.605 66.015 120.775 ;
        RECT 66.305 120.605 66.475 120.775 ;
        RECT 66.765 120.605 66.935 120.775 ;
        RECT 67.225 120.605 67.395 120.775 ;
        RECT 67.685 120.605 67.855 120.775 ;
        RECT 68.145 120.605 68.315 120.775 ;
        RECT 68.605 120.605 68.775 120.775 ;
        RECT 69.065 120.605 69.235 120.775 ;
        RECT 69.525 120.605 69.695 120.775 ;
        RECT 69.985 120.605 70.155 120.775 ;
        RECT 70.445 120.605 70.615 120.775 ;
        RECT 70.905 120.605 71.075 120.775 ;
        RECT 71.365 120.605 71.535 120.775 ;
        RECT 71.825 120.605 71.995 120.775 ;
        RECT 72.285 120.605 72.455 120.775 ;
        RECT 72.745 120.605 72.915 120.775 ;
        RECT 73.205 120.605 73.375 120.775 ;
        RECT 73.665 120.605 73.835 120.775 ;
        RECT 74.125 120.605 74.295 120.775 ;
        RECT 74.585 120.605 74.755 120.775 ;
        RECT 75.045 120.605 75.215 120.775 ;
        RECT 75.505 120.605 75.675 120.775 ;
        RECT 75.965 120.605 76.135 120.775 ;
        RECT 76.425 120.605 76.595 120.775 ;
        RECT 76.885 120.605 77.055 120.775 ;
        RECT 77.345 120.605 77.515 120.775 ;
        RECT 77.805 120.605 77.975 120.775 ;
        RECT 78.265 120.605 78.435 120.775 ;
        RECT 78.725 120.605 78.895 120.775 ;
        RECT 79.185 120.605 79.355 120.775 ;
        RECT 79.645 120.605 79.815 120.775 ;
        RECT 80.105 120.605 80.275 120.775 ;
        RECT 80.565 120.605 80.735 120.775 ;
        RECT 81.025 120.605 81.195 120.775 ;
        RECT 81.485 120.605 81.655 120.775 ;
        RECT 81.945 120.605 82.115 120.775 ;
        RECT 82.405 120.605 82.575 120.775 ;
        RECT 82.865 120.605 83.035 120.775 ;
        RECT 83.325 120.605 83.495 120.775 ;
        RECT 83.785 120.605 83.955 120.775 ;
        RECT 84.245 120.605 84.415 120.775 ;
        RECT 84.705 120.605 84.875 120.775 ;
        RECT 85.165 120.605 85.335 120.775 ;
        RECT 85.625 120.605 85.795 120.775 ;
        RECT 86.085 120.605 86.255 120.775 ;
        RECT 86.545 120.605 86.715 120.775 ;
        RECT 87.005 120.605 87.175 120.775 ;
        RECT 87.465 120.605 87.635 120.775 ;
        RECT 87.925 120.605 88.095 120.775 ;
        RECT 88.385 120.605 88.555 120.775 ;
        RECT 88.845 120.605 89.015 120.775 ;
        RECT 89.305 120.605 89.475 120.775 ;
        RECT 89.765 120.605 89.935 120.775 ;
        RECT 90.225 120.605 90.395 120.775 ;
        RECT 90.685 120.605 90.855 120.775 ;
        RECT 91.145 120.605 91.315 120.775 ;
        RECT 91.605 120.605 91.775 120.775 ;
        RECT 92.065 120.605 92.235 120.775 ;
        RECT 92.525 120.605 92.695 120.775 ;
        RECT 92.985 120.605 93.155 120.775 ;
        RECT 93.445 120.605 93.615 120.775 ;
        RECT 93.905 120.605 94.075 120.775 ;
        RECT 94.365 120.605 94.535 120.775 ;
        RECT 94.825 120.605 94.995 120.775 ;
        RECT 95.285 120.605 95.455 120.775 ;
        RECT 95.745 120.605 95.915 120.775 ;
        RECT 96.205 120.605 96.375 120.775 ;
        RECT 96.665 120.605 96.835 120.775 ;
        RECT 97.125 120.605 97.295 120.775 ;
        RECT 97.585 120.605 97.755 120.775 ;
        RECT 98.045 120.605 98.215 120.775 ;
        RECT 98.505 120.605 98.675 120.775 ;
        RECT 98.965 120.605 99.135 120.775 ;
        RECT 99.425 120.605 99.595 120.775 ;
        RECT 99.885 120.605 100.055 120.775 ;
        RECT 100.345 120.605 100.515 120.775 ;
        RECT 100.805 120.605 100.975 120.775 ;
        RECT 101.265 120.605 101.435 120.775 ;
        RECT 101.725 120.605 101.895 120.775 ;
        RECT 102.185 120.605 102.355 120.775 ;
        RECT 102.645 120.605 102.815 120.775 ;
        RECT 103.105 120.605 103.275 120.775 ;
        RECT 103.565 120.605 103.735 120.775 ;
        RECT 104.025 120.605 104.195 120.775 ;
        RECT 104.485 120.605 104.655 120.775 ;
        RECT 104.945 120.605 105.115 120.775 ;
        RECT 105.405 120.605 105.575 120.775 ;
        RECT 105.865 120.605 106.035 120.775 ;
        RECT 106.325 120.605 106.495 120.775 ;
        RECT 106.785 120.605 106.955 120.775 ;
        RECT 107.245 120.605 107.415 120.775 ;
        RECT 107.705 120.605 107.875 120.775 ;
        RECT 108.165 120.605 108.335 120.775 ;
        RECT 108.625 120.605 108.795 120.775 ;
        RECT 109.085 120.605 109.255 120.775 ;
        RECT 109.545 120.605 109.715 120.775 ;
        RECT 110.005 120.605 110.175 120.775 ;
        RECT 110.465 120.605 110.635 120.775 ;
        RECT 110.925 120.605 111.095 120.775 ;
        RECT 111.385 120.605 111.555 120.775 ;
        RECT 111.845 120.605 112.015 120.775 ;
        RECT 112.305 120.605 112.475 120.775 ;
        RECT 112.765 120.605 112.935 120.775 ;
        RECT 113.225 120.605 113.395 120.775 ;
        RECT 113.685 120.605 113.855 120.775 ;
        RECT 114.145 120.605 114.315 120.775 ;
        RECT 114.605 120.605 114.775 120.775 ;
        RECT 115.065 120.605 115.235 120.775 ;
        RECT 115.525 120.605 115.695 120.775 ;
        RECT 115.985 120.605 116.155 120.775 ;
        RECT 116.445 120.605 116.615 120.775 ;
        RECT 116.905 120.605 117.075 120.775 ;
        RECT 117.365 120.605 117.535 120.775 ;
        RECT 117.825 120.605 117.995 120.775 ;
        RECT 118.285 120.605 118.455 120.775 ;
        RECT 118.745 120.605 118.915 120.775 ;
        RECT 119.205 120.605 119.375 120.775 ;
        RECT 119.665 120.605 119.835 120.775 ;
        RECT 120.125 120.605 120.295 120.775 ;
        RECT 120.585 120.605 120.755 120.775 ;
        RECT 121.045 120.605 121.215 120.775 ;
        RECT 121.505 120.605 121.675 120.775 ;
        RECT 121.965 120.605 122.135 120.775 ;
        RECT 122.425 120.605 122.595 120.775 ;
        RECT 122.885 120.605 123.055 120.775 ;
        RECT 123.345 120.605 123.515 120.775 ;
        RECT 123.805 120.605 123.975 120.775 ;
        RECT 124.265 120.605 124.435 120.775 ;
        RECT 124.725 120.605 124.895 120.775 ;
        RECT 125.185 120.605 125.355 120.775 ;
        RECT 125.645 120.605 125.815 120.775 ;
        RECT 126.105 120.605 126.275 120.775 ;
        RECT 126.565 120.605 126.735 120.775 ;
        RECT 127.025 120.605 127.195 120.775 ;
        RECT 127.485 120.605 127.655 120.775 ;
        RECT 127.945 120.605 128.115 120.775 ;
        RECT 128.405 120.605 128.575 120.775 ;
        RECT 128.865 120.605 129.035 120.775 ;
        RECT 129.325 120.605 129.495 120.775 ;
        RECT 129.785 120.605 129.955 120.775 ;
        RECT 130.245 120.605 130.415 120.775 ;
        RECT 130.705 120.605 130.875 120.775 ;
        RECT 131.165 120.605 131.335 120.775 ;
        RECT 131.625 120.605 131.795 120.775 ;
        RECT 132.085 120.605 132.255 120.775 ;
        RECT 132.545 120.605 132.715 120.775 ;
        RECT 133.005 120.605 133.175 120.775 ;
        RECT 133.465 120.605 133.635 120.775 ;
        RECT 133.925 120.605 134.095 120.775 ;
        RECT 134.385 120.605 134.555 120.775 ;
        RECT 134.845 120.605 135.015 120.775 ;
        RECT 135.305 120.605 135.475 120.775 ;
        RECT 135.765 120.605 135.935 120.775 ;
        RECT 136.225 120.605 136.395 120.775 ;
        RECT 136.685 120.605 136.855 120.775 ;
        RECT 137.145 120.605 137.315 120.775 ;
        RECT 137.605 120.605 137.775 120.775 ;
        RECT 138.065 120.605 138.235 120.775 ;
        RECT 138.525 120.605 138.695 120.775 ;
        RECT 138.985 120.605 139.155 120.775 ;
        RECT 50.665 117.885 50.835 118.055 ;
        RECT 51.125 117.885 51.295 118.055 ;
        RECT 51.585 117.885 51.755 118.055 ;
        RECT 52.045 117.885 52.215 118.055 ;
        RECT 52.505 117.885 52.675 118.055 ;
        RECT 52.965 117.885 53.135 118.055 ;
        RECT 53.425 117.885 53.595 118.055 ;
        RECT 53.885 117.885 54.055 118.055 ;
        RECT 54.345 117.885 54.515 118.055 ;
        RECT 54.805 117.885 54.975 118.055 ;
        RECT 55.265 117.885 55.435 118.055 ;
        RECT 55.725 117.885 55.895 118.055 ;
        RECT 56.185 117.885 56.355 118.055 ;
        RECT 56.645 117.885 56.815 118.055 ;
        RECT 57.105 117.885 57.275 118.055 ;
        RECT 57.565 117.885 57.735 118.055 ;
        RECT 58.025 117.885 58.195 118.055 ;
        RECT 58.485 117.885 58.655 118.055 ;
        RECT 58.945 117.885 59.115 118.055 ;
        RECT 59.405 117.885 59.575 118.055 ;
        RECT 59.865 117.885 60.035 118.055 ;
        RECT 60.325 117.885 60.495 118.055 ;
        RECT 60.785 117.885 60.955 118.055 ;
        RECT 61.245 117.885 61.415 118.055 ;
        RECT 61.705 117.885 61.875 118.055 ;
        RECT 62.165 117.885 62.335 118.055 ;
        RECT 62.625 117.885 62.795 118.055 ;
        RECT 63.085 117.885 63.255 118.055 ;
        RECT 63.545 117.885 63.715 118.055 ;
        RECT 64.005 117.885 64.175 118.055 ;
        RECT 64.465 117.885 64.635 118.055 ;
        RECT 64.925 117.885 65.095 118.055 ;
        RECT 65.385 117.885 65.555 118.055 ;
        RECT 65.845 117.885 66.015 118.055 ;
        RECT 66.305 117.885 66.475 118.055 ;
        RECT 66.765 117.885 66.935 118.055 ;
        RECT 67.225 117.885 67.395 118.055 ;
        RECT 67.685 117.885 67.855 118.055 ;
        RECT 68.145 117.885 68.315 118.055 ;
        RECT 68.605 117.885 68.775 118.055 ;
        RECT 69.065 117.885 69.235 118.055 ;
        RECT 69.525 117.885 69.695 118.055 ;
        RECT 69.985 117.885 70.155 118.055 ;
        RECT 70.445 117.885 70.615 118.055 ;
        RECT 70.905 117.885 71.075 118.055 ;
        RECT 71.365 117.885 71.535 118.055 ;
        RECT 71.825 117.885 71.995 118.055 ;
        RECT 72.285 117.885 72.455 118.055 ;
        RECT 72.745 117.885 72.915 118.055 ;
        RECT 73.205 117.885 73.375 118.055 ;
        RECT 73.665 117.885 73.835 118.055 ;
        RECT 74.125 117.885 74.295 118.055 ;
        RECT 74.585 117.885 74.755 118.055 ;
        RECT 75.045 117.885 75.215 118.055 ;
        RECT 75.505 117.885 75.675 118.055 ;
        RECT 75.965 117.885 76.135 118.055 ;
        RECT 76.425 117.885 76.595 118.055 ;
        RECT 76.885 117.885 77.055 118.055 ;
        RECT 77.345 117.885 77.515 118.055 ;
        RECT 77.805 117.885 77.975 118.055 ;
        RECT 78.265 117.885 78.435 118.055 ;
        RECT 78.725 117.885 78.895 118.055 ;
        RECT 79.185 117.885 79.355 118.055 ;
        RECT 79.645 117.885 79.815 118.055 ;
        RECT 80.105 117.885 80.275 118.055 ;
        RECT 80.565 117.885 80.735 118.055 ;
        RECT 81.025 117.885 81.195 118.055 ;
        RECT 81.485 117.885 81.655 118.055 ;
        RECT 81.945 117.885 82.115 118.055 ;
        RECT 82.405 117.885 82.575 118.055 ;
        RECT 82.865 117.885 83.035 118.055 ;
        RECT 83.325 117.885 83.495 118.055 ;
        RECT 83.785 117.885 83.955 118.055 ;
        RECT 84.245 117.885 84.415 118.055 ;
        RECT 84.705 117.885 84.875 118.055 ;
        RECT 85.165 117.885 85.335 118.055 ;
        RECT 85.625 117.885 85.795 118.055 ;
        RECT 86.085 117.885 86.255 118.055 ;
        RECT 86.545 117.885 86.715 118.055 ;
        RECT 87.005 117.885 87.175 118.055 ;
        RECT 87.465 117.885 87.635 118.055 ;
        RECT 87.925 117.885 88.095 118.055 ;
        RECT 88.385 117.885 88.555 118.055 ;
        RECT 88.845 117.885 89.015 118.055 ;
        RECT 89.305 117.885 89.475 118.055 ;
        RECT 89.765 117.885 89.935 118.055 ;
        RECT 90.225 117.885 90.395 118.055 ;
        RECT 90.685 117.885 90.855 118.055 ;
        RECT 91.145 117.885 91.315 118.055 ;
        RECT 91.605 117.885 91.775 118.055 ;
        RECT 92.065 117.885 92.235 118.055 ;
        RECT 92.525 117.885 92.695 118.055 ;
        RECT 92.985 117.885 93.155 118.055 ;
        RECT 93.445 117.885 93.615 118.055 ;
        RECT 93.905 117.885 94.075 118.055 ;
        RECT 94.365 117.885 94.535 118.055 ;
        RECT 94.825 117.885 94.995 118.055 ;
        RECT 95.285 117.885 95.455 118.055 ;
        RECT 95.745 117.885 95.915 118.055 ;
        RECT 96.205 117.885 96.375 118.055 ;
        RECT 96.665 117.885 96.835 118.055 ;
        RECT 97.125 117.885 97.295 118.055 ;
        RECT 97.585 117.885 97.755 118.055 ;
        RECT 98.045 117.885 98.215 118.055 ;
        RECT 98.505 117.885 98.675 118.055 ;
        RECT 98.965 117.885 99.135 118.055 ;
        RECT 99.425 117.885 99.595 118.055 ;
        RECT 99.885 117.885 100.055 118.055 ;
        RECT 100.345 117.885 100.515 118.055 ;
        RECT 100.805 117.885 100.975 118.055 ;
        RECT 101.265 117.885 101.435 118.055 ;
        RECT 101.725 117.885 101.895 118.055 ;
        RECT 102.185 117.885 102.355 118.055 ;
        RECT 102.645 117.885 102.815 118.055 ;
        RECT 103.105 117.885 103.275 118.055 ;
        RECT 103.565 117.885 103.735 118.055 ;
        RECT 104.025 117.885 104.195 118.055 ;
        RECT 104.485 117.885 104.655 118.055 ;
        RECT 104.945 117.885 105.115 118.055 ;
        RECT 105.405 117.885 105.575 118.055 ;
        RECT 105.865 117.885 106.035 118.055 ;
        RECT 106.325 117.885 106.495 118.055 ;
        RECT 106.785 117.885 106.955 118.055 ;
        RECT 107.245 117.885 107.415 118.055 ;
        RECT 107.705 117.885 107.875 118.055 ;
        RECT 108.165 117.885 108.335 118.055 ;
        RECT 108.625 117.885 108.795 118.055 ;
        RECT 109.085 117.885 109.255 118.055 ;
        RECT 109.545 117.885 109.715 118.055 ;
        RECT 110.005 117.885 110.175 118.055 ;
        RECT 110.465 117.885 110.635 118.055 ;
        RECT 110.925 117.885 111.095 118.055 ;
        RECT 111.385 117.885 111.555 118.055 ;
        RECT 111.845 117.885 112.015 118.055 ;
        RECT 112.305 117.885 112.475 118.055 ;
        RECT 112.765 117.885 112.935 118.055 ;
        RECT 113.225 117.885 113.395 118.055 ;
        RECT 113.685 117.885 113.855 118.055 ;
        RECT 114.145 117.885 114.315 118.055 ;
        RECT 114.605 117.885 114.775 118.055 ;
        RECT 115.065 117.885 115.235 118.055 ;
        RECT 115.525 117.885 115.695 118.055 ;
        RECT 115.985 117.885 116.155 118.055 ;
        RECT 116.445 117.885 116.615 118.055 ;
        RECT 116.905 117.885 117.075 118.055 ;
        RECT 117.365 117.885 117.535 118.055 ;
        RECT 117.825 117.885 117.995 118.055 ;
        RECT 118.285 117.885 118.455 118.055 ;
        RECT 118.745 117.885 118.915 118.055 ;
        RECT 119.205 117.885 119.375 118.055 ;
        RECT 119.665 117.885 119.835 118.055 ;
        RECT 120.125 117.885 120.295 118.055 ;
        RECT 120.585 117.885 120.755 118.055 ;
        RECT 121.045 117.885 121.215 118.055 ;
        RECT 121.505 117.885 121.675 118.055 ;
        RECT 121.965 117.885 122.135 118.055 ;
        RECT 122.425 117.885 122.595 118.055 ;
        RECT 122.885 117.885 123.055 118.055 ;
        RECT 123.345 117.885 123.515 118.055 ;
        RECT 123.805 117.885 123.975 118.055 ;
        RECT 124.265 117.885 124.435 118.055 ;
        RECT 124.725 117.885 124.895 118.055 ;
        RECT 125.185 117.885 125.355 118.055 ;
        RECT 125.645 117.885 125.815 118.055 ;
        RECT 126.105 117.885 126.275 118.055 ;
        RECT 126.565 117.885 126.735 118.055 ;
        RECT 127.025 117.885 127.195 118.055 ;
        RECT 127.485 117.885 127.655 118.055 ;
        RECT 127.945 117.885 128.115 118.055 ;
        RECT 128.405 117.885 128.575 118.055 ;
        RECT 128.865 117.885 129.035 118.055 ;
        RECT 129.325 117.885 129.495 118.055 ;
        RECT 129.785 117.885 129.955 118.055 ;
        RECT 130.245 117.885 130.415 118.055 ;
        RECT 130.705 117.885 130.875 118.055 ;
        RECT 131.165 117.885 131.335 118.055 ;
        RECT 131.625 117.885 131.795 118.055 ;
        RECT 132.085 117.885 132.255 118.055 ;
        RECT 132.545 117.885 132.715 118.055 ;
        RECT 133.005 117.885 133.175 118.055 ;
        RECT 133.465 117.885 133.635 118.055 ;
        RECT 133.925 117.885 134.095 118.055 ;
        RECT 134.385 117.885 134.555 118.055 ;
        RECT 134.845 117.885 135.015 118.055 ;
        RECT 135.305 117.885 135.475 118.055 ;
        RECT 135.765 117.885 135.935 118.055 ;
        RECT 136.225 117.885 136.395 118.055 ;
        RECT 136.685 117.885 136.855 118.055 ;
        RECT 137.145 117.885 137.315 118.055 ;
        RECT 137.605 117.885 137.775 118.055 ;
        RECT 138.065 117.885 138.235 118.055 ;
        RECT 138.525 117.885 138.695 118.055 ;
        RECT 138.985 117.885 139.155 118.055 ;
        RECT 50.665 115.165 50.835 115.335 ;
        RECT 51.125 115.165 51.295 115.335 ;
        RECT 51.585 115.165 51.755 115.335 ;
        RECT 52.045 115.165 52.215 115.335 ;
        RECT 52.505 115.165 52.675 115.335 ;
        RECT 52.965 115.165 53.135 115.335 ;
        RECT 53.425 115.165 53.595 115.335 ;
        RECT 53.885 115.165 54.055 115.335 ;
        RECT 54.345 115.165 54.515 115.335 ;
        RECT 54.805 115.165 54.975 115.335 ;
        RECT 55.265 115.165 55.435 115.335 ;
        RECT 55.725 115.165 55.895 115.335 ;
        RECT 56.185 115.165 56.355 115.335 ;
        RECT 56.645 115.165 56.815 115.335 ;
        RECT 57.105 115.165 57.275 115.335 ;
        RECT 57.565 115.165 57.735 115.335 ;
        RECT 58.025 115.165 58.195 115.335 ;
        RECT 58.485 115.165 58.655 115.335 ;
        RECT 58.945 115.165 59.115 115.335 ;
        RECT 59.405 115.165 59.575 115.335 ;
        RECT 59.865 115.165 60.035 115.335 ;
        RECT 60.325 115.165 60.495 115.335 ;
        RECT 60.785 115.165 60.955 115.335 ;
        RECT 61.245 115.165 61.415 115.335 ;
        RECT 61.705 115.165 61.875 115.335 ;
        RECT 62.165 115.165 62.335 115.335 ;
        RECT 62.625 115.165 62.795 115.335 ;
        RECT 63.085 115.165 63.255 115.335 ;
        RECT 63.545 115.165 63.715 115.335 ;
        RECT 64.005 115.165 64.175 115.335 ;
        RECT 64.465 115.165 64.635 115.335 ;
        RECT 64.925 115.165 65.095 115.335 ;
        RECT 65.385 115.165 65.555 115.335 ;
        RECT 65.845 115.165 66.015 115.335 ;
        RECT 66.305 115.165 66.475 115.335 ;
        RECT 66.765 115.165 66.935 115.335 ;
        RECT 67.225 115.165 67.395 115.335 ;
        RECT 67.685 115.165 67.855 115.335 ;
        RECT 68.145 115.165 68.315 115.335 ;
        RECT 68.605 115.165 68.775 115.335 ;
        RECT 69.065 115.165 69.235 115.335 ;
        RECT 69.525 115.165 69.695 115.335 ;
        RECT 69.985 115.165 70.155 115.335 ;
        RECT 70.445 115.165 70.615 115.335 ;
        RECT 70.905 115.165 71.075 115.335 ;
        RECT 71.365 115.165 71.535 115.335 ;
        RECT 71.825 115.165 71.995 115.335 ;
        RECT 72.285 115.165 72.455 115.335 ;
        RECT 72.745 115.165 72.915 115.335 ;
        RECT 73.205 115.165 73.375 115.335 ;
        RECT 73.665 115.165 73.835 115.335 ;
        RECT 74.125 115.165 74.295 115.335 ;
        RECT 74.585 115.165 74.755 115.335 ;
        RECT 75.045 115.165 75.215 115.335 ;
        RECT 75.505 115.165 75.675 115.335 ;
        RECT 75.965 115.165 76.135 115.335 ;
        RECT 76.425 115.165 76.595 115.335 ;
        RECT 76.885 115.165 77.055 115.335 ;
        RECT 77.345 115.165 77.515 115.335 ;
        RECT 77.805 115.165 77.975 115.335 ;
        RECT 78.265 115.165 78.435 115.335 ;
        RECT 78.725 115.165 78.895 115.335 ;
        RECT 79.185 115.165 79.355 115.335 ;
        RECT 79.645 115.165 79.815 115.335 ;
        RECT 80.105 115.165 80.275 115.335 ;
        RECT 80.565 115.165 80.735 115.335 ;
        RECT 81.025 115.165 81.195 115.335 ;
        RECT 81.485 115.165 81.655 115.335 ;
        RECT 81.945 115.165 82.115 115.335 ;
        RECT 82.405 115.165 82.575 115.335 ;
        RECT 82.865 115.165 83.035 115.335 ;
        RECT 83.325 115.165 83.495 115.335 ;
        RECT 83.785 115.165 83.955 115.335 ;
        RECT 84.245 115.165 84.415 115.335 ;
        RECT 84.705 115.165 84.875 115.335 ;
        RECT 85.165 115.165 85.335 115.335 ;
        RECT 85.625 115.165 85.795 115.335 ;
        RECT 86.085 115.165 86.255 115.335 ;
        RECT 86.545 115.165 86.715 115.335 ;
        RECT 87.005 115.165 87.175 115.335 ;
        RECT 87.465 115.165 87.635 115.335 ;
        RECT 87.925 115.165 88.095 115.335 ;
        RECT 88.385 115.165 88.555 115.335 ;
        RECT 88.845 115.165 89.015 115.335 ;
        RECT 89.305 115.165 89.475 115.335 ;
        RECT 89.765 115.165 89.935 115.335 ;
        RECT 90.225 115.165 90.395 115.335 ;
        RECT 90.685 115.165 90.855 115.335 ;
        RECT 91.145 115.165 91.315 115.335 ;
        RECT 91.605 115.165 91.775 115.335 ;
        RECT 92.065 115.165 92.235 115.335 ;
        RECT 92.525 115.165 92.695 115.335 ;
        RECT 92.985 115.165 93.155 115.335 ;
        RECT 93.445 115.165 93.615 115.335 ;
        RECT 93.905 115.165 94.075 115.335 ;
        RECT 94.365 115.165 94.535 115.335 ;
        RECT 94.825 115.165 94.995 115.335 ;
        RECT 95.285 115.165 95.455 115.335 ;
        RECT 95.745 115.165 95.915 115.335 ;
        RECT 96.205 115.165 96.375 115.335 ;
        RECT 96.665 115.165 96.835 115.335 ;
        RECT 97.125 115.165 97.295 115.335 ;
        RECT 97.585 115.165 97.755 115.335 ;
        RECT 98.045 115.165 98.215 115.335 ;
        RECT 98.505 115.165 98.675 115.335 ;
        RECT 98.965 115.165 99.135 115.335 ;
        RECT 99.425 115.165 99.595 115.335 ;
        RECT 99.885 115.165 100.055 115.335 ;
        RECT 100.345 115.165 100.515 115.335 ;
        RECT 100.805 115.165 100.975 115.335 ;
        RECT 101.265 115.165 101.435 115.335 ;
        RECT 101.725 115.165 101.895 115.335 ;
        RECT 102.185 115.165 102.355 115.335 ;
        RECT 102.645 115.165 102.815 115.335 ;
        RECT 103.105 115.165 103.275 115.335 ;
        RECT 103.565 115.165 103.735 115.335 ;
        RECT 104.025 115.165 104.195 115.335 ;
        RECT 104.485 115.165 104.655 115.335 ;
        RECT 104.945 115.165 105.115 115.335 ;
        RECT 105.405 115.165 105.575 115.335 ;
        RECT 105.865 115.165 106.035 115.335 ;
        RECT 106.325 115.165 106.495 115.335 ;
        RECT 106.785 115.165 106.955 115.335 ;
        RECT 107.245 115.165 107.415 115.335 ;
        RECT 107.705 115.165 107.875 115.335 ;
        RECT 108.165 115.165 108.335 115.335 ;
        RECT 108.625 115.165 108.795 115.335 ;
        RECT 109.085 115.165 109.255 115.335 ;
        RECT 109.545 115.165 109.715 115.335 ;
        RECT 110.005 115.165 110.175 115.335 ;
        RECT 110.465 115.165 110.635 115.335 ;
        RECT 110.925 115.165 111.095 115.335 ;
        RECT 111.385 115.165 111.555 115.335 ;
        RECT 111.845 115.165 112.015 115.335 ;
        RECT 112.305 115.165 112.475 115.335 ;
        RECT 112.765 115.165 112.935 115.335 ;
        RECT 113.225 115.165 113.395 115.335 ;
        RECT 113.685 115.165 113.855 115.335 ;
        RECT 114.145 115.165 114.315 115.335 ;
        RECT 114.605 115.165 114.775 115.335 ;
        RECT 115.065 115.165 115.235 115.335 ;
        RECT 115.525 115.165 115.695 115.335 ;
        RECT 115.985 115.165 116.155 115.335 ;
        RECT 116.445 115.165 116.615 115.335 ;
        RECT 116.905 115.165 117.075 115.335 ;
        RECT 117.365 115.165 117.535 115.335 ;
        RECT 117.825 115.165 117.995 115.335 ;
        RECT 118.285 115.165 118.455 115.335 ;
        RECT 118.745 115.165 118.915 115.335 ;
        RECT 119.205 115.165 119.375 115.335 ;
        RECT 119.665 115.165 119.835 115.335 ;
        RECT 120.125 115.165 120.295 115.335 ;
        RECT 120.585 115.165 120.755 115.335 ;
        RECT 121.045 115.165 121.215 115.335 ;
        RECT 121.505 115.165 121.675 115.335 ;
        RECT 121.965 115.165 122.135 115.335 ;
        RECT 122.425 115.165 122.595 115.335 ;
        RECT 122.885 115.165 123.055 115.335 ;
        RECT 123.345 115.165 123.515 115.335 ;
        RECT 123.805 115.165 123.975 115.335 ;
        RECT 124.265 115.165 124.435 115.335 ;
        RECT 124.725 115.165 124.895 115.335 ;
        RECT 125.185 115.165 125.355 115.335 ;
        RECT 125.645 115.165 125.815 115.335 ;
        RECT 126.105 115.165 126.275 115.335 ;
        RECT 126.565 115.165 126.735 115.335 ;
        RECT 127.025 115.165 127.195 115.335 ;
        RECT 127.485 115.165 127.655 115.335 ;
        RECT 127.945 115.165 128.115 115.335 ;
        RECT 128.405 115.165 128.575 115.335 ;
        RECT 128.865 115.165 129.035 115.335 ;
        RECT 129.325 115.165 129.495 115.335 ;
        RECT 129.785 115.165 129.955 115.335 ;
        RECT 130.245 115.165 130.415 115.335 ;
        RECT 130.705 115.165 130.875 115.335 ;
        RECT 131.165 115.165 131.335 115.335 ;
        RECT 131.625 115.165 131.795 115.335 ;
        RECT 132.085 115.165 132.255 115.335 ;
        RECT 132.545 115.165 132.715 115.335 ;
        RECT 133.005 115.165 133.175 115.335 ;
        RECT 133.465 115.165 133.635 115.335 ;
        RECT 133.925 115.165 134.095 115.335 ;
        RECT 134.385 115.165 134.555 115.335 ;
        RECT 134.845 115.165 135.015 115.335 ;
        RECT 135.305 115.165 135.475 115.335 ;
        RECT 135.765 115.165 135.935 115.335 ;
        RECT 136.225 115.165 136.395 115.335 ;
        RECT 136.685 115.165 136.855 115.335 ;
        RECT 137.145 115.165 137.315 115.335 ;
        RECT 137.605 115.165 137.775 115.335 ;
        RECT 138.065 115.165 138.235 115.335 ;
        RECT 138.525 115.165 138.695 115.335 ;
        RECT 138.985 115.165 139.155 115.335 ;
        RECT 50.665 112.445 50.835 112.615 ;
        RECT 51.125 112.445 51.295 112.615 ;
        RECT 51.585 112.445 51.755 112.615 ;
        RECT 52.045 112.445 52.215 112.615 ;
        RECT 52.505 112.445 52.675 112.615 ;
        RECT 52.965 112.445 53.135 112.615 ;
        RECT 53.425 112.445 53.595 112.615 ;
        RECT 53.885 112.445 54.055 112.615 ;
        RECT 54.345 112.445 54.515 112.615 ;
        RECT 54.805 112.445 54.975 112.615 ;
        RECT 55.265 112.445 55.435 112.615 ;
        RECT 55.725 112.445 55.895 112.615 ;
        RECT 56.185 112.445 56.355 112.615 ;
        RECT 56.645 112.445 56.815 112.615 ;
        RECT 57.105 112.445 57.275 112.615 ;
        RECT 57.565 112.445 57.735 112.615 ;
        RECT 58.025 112.445 58.195 112.615 ;
        RECT 58.485 112.445 58.655 112.615 ;
        RECT 58.945 112.445 59.115 112.615 ;
        RECT 59.405 112.445 59.575 112.615 ;
        RECT 59.865 112.445 60.035 112.615 ;
        RECT 60.325 112.445 60.495 112.615 ;
        RECT 60.785 112.445 60.955 112.615 ;
        RECT 61.245 112.445 61.415 112.615 ;
        RECT 61.705 112.445 61.875 112.615 ;
        RECT 62.165 112.445 62.335 112.615 ;
        RECT 62.625 112.445 62.795 112.615 ;
        RECT 63.085 112.445 63.255 112.615 ;
        RECT 63.545 112.445 63.715 112.615 ;
        RECT 64.005 112.445 64.175 112.615 ;
        RECT 64.465 112.445 64.635 112.615 ;
        RECT 64.925 112.445 65.095 112.615 ;
        RECT 65.385 112.445 65.555 112.615 ;
        RECT 65.845 112.445 66.015 112.615 ;
        RECT 66.305 112.445 66.475 112.615 ;
        RECT 66.765 112.445 66.935 112.615 ;
        RECT 67.225 112.445 67.395 112.615 ;
        RECT 67.685 112.445 67.855 112.615 ;
        RECT 68.145 112.445 68.315 112.615 ;
        RECT 68.605 112.445 68.775 112.615 ;
        RECT 69.065 112.445 69.235 112.615 ;
        RECT 69.525 112.445 69.695 112.615 ;
        RECT 69.985 112.445 70.155 112.615 ;
        RECT 70.445 112.445 70.615 112.615 ;
        RECT 70.905 112.445 71.075 112.615 ;
        RECT 71.365 112.445 71.535 112.615 ;
        RECT 71.825 112.445 71.995 112.615 ;
        RECT 72.285 112.445 72.455 112.615 ;
        RECT 72.745 112.445 72.915 112.615 ;
        RECT 73.205 112.445 73.375 112.615 ;
        RECT 73.665 112.445 73.835 112.615 ;
        RECT 74.125 112.445 74.295 112.615 ;
        RECT 74.585 112.445 74.755 112.615 ;
        RECT 75.045 112.445 75.215 112.615 ;
        RECT 75.505 112.445 75.675 112.615 ;
        RECT 75.965 112.445 76.135 112.615 ;
        RECT 76.425 112.445 76.595 112.615 ;
        RECT 76.885 112.445 77.055 112.615 ;
        RECT 77.345 112.445 77.515 112.615 ;
        RECT 77.805 112.445 77.975 112.615 ;
        RECT 78.265 112.445 78.435 112.615 ;
        RECT 78.725 112.445 78.895 112.615 ;
        RECT 79.185 112.445 79.355 112.615 ;
        RECT 79.645 112.445 79.815 112.615 ;
        RECT 80.105 112.445 80.275 112.615 ;
        RECT 80.565 112.445 80.735 112.615 ;
        RECT 81.025 112.445 81.195 112.615 ;
        RECT 81.485 112.445 81.655 112.615 ;
        RECT 81.945 112.445 82.115 112.615 ;
        RECT 82.405 112.445 82.575 112.615 ;
        RECT 82.865 112.445 83.035 112.615 ;
        RECT 83.325 112.445 83.495 112.615 ;
        RECT 83.785 112.445 83.955 112.615 ;
        RECT 84.245 112.445 84.415 112.615 ;
        RECT 84.705 112.445 84.875 112.615 ;
        RECT 85.165 112.445 85.335 112.615 ;
        RECT 85.625 112.445 85.795 112.615 ;
        RECT 86.085 112.445 86.255 112.615 ;
        RECT 86.545 112.445 86.715 112.615 ;
        RECT 87.005 112.445 87.175 112.615 ;
        RECT 87.465 112.445 87.635 112.615 ;
        RECT 87.925 112.445 88.095 112.615 ;
        RECT 88.385 112.445 88.555 112.615 ;
        RECT 88.845 112.445 89.015 112.615 ;
        RECT 89.305 112.445 89.475 112.615 ;
        RECT 89.765 112.445 89.935 112.615 ;
        RECT 90.225 112.445 90.395 112.615 ;
        RECT 90.685 112.445 90.855 112.615 ;
        RECT 91.145 112.445 91.315 112.615 ;
        RECT 91.605 112.445 91.775 112.615 ;
        RECT 92.065 112.445 92.235 112.615 ;
        RECT 92.525 112.445 92.695 112.615 ;
        RECT 92.985 112.445 93.155 112.615 ;
        RECT 93.445 112.445 93.615 112.615 ;
        RECT 93.905 112.445 94.075 112.615 ;
        RECT 94.365 112.445 94.535 112.615 ;
        RECT 94.825 112.445 94.995 112.615 ;
        RECT 95.285 112.445 95.455 112.615 ;
        RECT 95.745 112.445 95.915 112.615 ;
        RECT 96.205 112.445 96.375 112.615 ;
        RECT 96.665 112.445 96.835 112.615 ;
        RECT 97.125 112.445 97.295 112.615 ;
        RECT 97.585 112.445 97.755 112.615 ;
        RECT 98.045 112.445 98.215 112.615 ;
        RECT 98.505 112.445 98.675 112.615 ;
        RECT 98.965 112.445 99.135 112.615 ;
        RECT 99.425 112.445 99.595 112.615 ;
        RECT 99.885 112.445 100.055 112.615 ;
        RECT 100.345 112.445 100.515 112.615 ;
        RECT 100.805 112.445 100.975 112.615 ;
        RECT 101.265 112.445 101.435 112.615 ;
        RECT 101.725 112.445 101.895 112.615 ;
        RECT 102.185 112.445 102.355 112.615 ;
        RECT 102.645 112.445 102.815 112.615 ;
        RECT 103.105 112.445 103.275 112.615 ;
        RECT 103.565 112.445 103.735 112.615 ;
        RECT 104.025 112.445 104.195 112.615 ;
        RECT 104.485 112.445 104.655 112.615 ;
        RECT 104.945 112.445 105.115 112.615 ;
        RECT 105.405 112.445 105.575 112.615 ;
        RECT 105.865 112.445 106.035 112.615 ;
        RECT 106.325 112.445 106.495 112.615 ;
        RECT 106.785 112.445 106.955 112.615 ;
        RECT 107.245 112.445 107.415 112.615 ;
        RECT 107.705 112.445 107.875 112.615 ;
        RECT 108.165 112.445 108.335 112.615 ;
        RECT 108.625 112.445 108.795 112.615 ;
        RECT 109.085 112.445 109.255 112.615 ;
        RECT 109.545 112.445 109.715 112.615 ;
        RECT 110.005 112.445 110.175 112.615 ;
        RECT 110.465 112.445 110.635 112.615 ;
        RECT 110.925 112.445 111.095 112.615 ;
        RECT 111.385 112.445 111.555 112.615 ;
        RECT 111.845 112.445 112.015 112.615 ;
        RECT 112.305 112.445 112.475 112.615 ;
        RECT 112.765 112.445 112.935 112.615 ;
        RECT 113.225 112.445 113.395 112.615 ;
        RECT 113.685 112.445 113.855 112.615 ;
        RECT 114.145 112.445 114.315 112.615 ;
        RECT 114.605 112.445 114.775 112.615 ;
        RECT 115.065 112.445 115.235 112.615 ;
        RECT 115.525 112.445 115.695 112.615 ;
        RECT 115.985 112.445 116.155 112.615 ;
        RECT 116.445 112.445 116.615 112.615 ;
        RECT 116.905 112.445 117.075 112.615 ;
        RECT 117.365 112.445 117.535 112.615 ;
        RECT 117.825 112.445 117.995 112.615 ;
        RECT 118.285 112.445 118.455 112.615 ;
        RECT 118.745 112.445 118.915 112.615 ;
        RECT 119.205 112.445 119.375 112.615 ;
        RECT 119.665 112.445 119.835 112.615 ;
        RECT 120.125 112.445 120.295 112.615 ;
        RECT 120.585 112.445 120.755 112.615 ;
        RECT 121.045 112.445 121.215 112.615 ;
        RECT 121.505 112.445 121.675 112.615 ;
        RECT 121.965 112.445 122.135 112.615 ;
        RECT 122.425 112.445 122.595 112.615 ;
        RECT 122.885 112.445 123.055 112.615 ;
        RECT 123.345 112.445 123.515 112.615 ;
        RECT 123.805 112.445 123.975 112.615 ;
        RECT 124.265 112.445 124.435 112.615 ;
        RECT 124.725 112.445 124.895 112.615 ;
        RECT 125.185 112.445 125.355 112.615 ;
        RECT 125.645 112.445 125.815 112.615 ;
        RECT 126.105 112.445 126.275 112.615 ;
        RECT 126.565 112.445 126.735 112.615 ;
        RECT 127.025 112.445 127.195 112.615 ;
        RECT 127.485 112.445 127.655 112.615 ;
        RECT 127.945 112.445 128.115 112.615 ;
        RECT 128.405 112.445 128.575 112.615 ;
        RECT 128.865 112.445 129.035 112.615 ;
        RECT 129.325 112.445 129.495 112.615 ;
        RECT 129.785 112.445 129.955 112.615 ;
        RECT 130.245 112.445 130.415 112.615 ;
        RECT 130.705 112.445 130.875 112.615 ;
        RECT 131.165 112.445 131.335 112.615 ;
        RECT 131.625 112.445 131.795 112.615 ;
        RECT 132.085 112.445 132.255 112.615 ;
        RECT 132.545 112.445 132.715 112.615 ;
        RECT 133.005 112.445 133.175 112.615 ;
        RECT 133.465 112.445 133.635 112.615 ;
        RECT 133.925 112.445 134.095 112.615 ;
        RECT 134.385 112.445 134.555 112.615 ;
        RECT 134.845 112.445 135.015 112.615 ;
        RECT 135.305 112.445 135.475 112.615 ;
        RECT 135.765 112.445 135.935 112.615 ;
        RECT 136.225 112.445 136.395 112.615 ;
        RECT 136.685 112.445 136.855 112.615 ;
        RECT 137.145 112.445 137.315 112.615 ;
        RECT 137.605 112.445 137.775 112.615 ;
        RECT 138.065 112.445 138.235 112.615 ;
        RECT 138.525 112.445 138.695 112.615 ;
        RECT 138.985 112.445 139.155 112.615 ;
        RECT 50.665 109.725 50.835 109.895 ;
        RECT 51.125 109.725 51.295 109.895 ;
        RECT 51.585 109.725 51.755 109.895 ;
        RECT 52.045 109.725 52.215 109.895 ;
        RECT 52.505 109.725 52.675 109.895 ;
        RECT 52.965 109.725 53.135 109.895 ;
        RECT 53.425 109.725 53.595 109.895 ;
        RECT 53.885 109.725 54.055 109.895 ;
        RECT 54.345 109.725 54.515 109.895 ;
        RECT 54.805 109.725 54.975 109.895 ;
        RECT 55.265 109.725 55.435 109.895 ;
        RECT 55.725 109.725 55.895 109.895 ;
        RECT 56.185 109.725 56.355 109.895 ;
        RECT 56.645 109.725 56.815 109.895 ;
        RECT 57.105 109.725 57.275 109.895 ;
        RECT 57.565 109.725 57.735 109.895 ;
        RECT 58.025 109.725 58.195 109.895 ;
        RECT 58.485 109.725 58.655 109.895 ;
        RECT 58.945 109.725 59.115 109.895 ;
        RECT 59.405 109.725 59.575 109.895 ;
        RECT 59.865 109.725 60.035 109.895 ;
        RECT 60.325 109.725 60.495 109.895 ;
        RECT 60.785 109.725 60.955 109.895 ;
        RECT 61.245 109.725 61.415 109.895 ;
        RECT 61.705 109.725 61.875 109.895 ;
        RECT 62.165 109.725 62.335 109.895 ;
        RECT 62.625 109.725 62.795 109.895 ;
        RECT 63.085 109.725 63.255 109.895 ;
        RECT 63.545 109.725 63.715 109.895 ;
        RECT 64.005 109.725 64.175 109.895 ;
        RECT 64.465 109.725 64.635 109.895 ;
        RECT 64.925 109.725 65.095 109.895 ;
        RECT 65.385 109.725 65.555 109.895 ;
        RECT 65.845 109.725 66.015 109.895 ;
        RECT 66.305 109.725 66.475 109.895 ;
        RECT 66.765 109.725 66.935 109.895 ;
        RECT 67.225 109.725 67.395 109.895 ;
        RECT 67.685 109.725 67.855 109.895 ;
        RECT 68.145 109.725 68.315 109.895 ;
        RECT 68.605 109.725 68.775 109.895 ;
        RECT 69.065 109.725 69.235 109.895 ;
        RECT 69.525 109.725 69.695 109.895 ;
        RECT 69.985 109.725 70.155 109.895 ;
        RECT 70.445 109.725 70.615 109.895 ;
        RECT 70.905 109.725 71.075 109.895 ;
        RECT 71.365 109.725 71.535 109.895 ;
        RECT 71.825 109.725 71.995 109.895 ;
        RECT 72.285 109.725 72.455 109.895 ;
        RECT 72.745 109.725 72.915 109.895 ;
        RECT 73.205 109.725 73.375 109.895 ;
        RECT 73.665 109.725 73.835 109.895 ;
        RECT 74.125 109.725 74.295 109.895 ;
        RECT 74.585 109.725 74.755 109.895 ;
        RECT 75.045 109.725 75.215 109.895 ;
        RECT 75.505 109.725 75.675 109.895 ;
        RECT 75.965 109.725 76.135 109.895 ;
        RECT 76.425 109.725 76.595 109.895 ;
        RECT 76.885 109.725 77.055 109.895 ;
        RECT 77.345 109.725 77.515 109.895 ;
        RECT 77.805 109.725 77.975 109.895 ;
        RECT 78.265 109.725 78.435 109.895 ;
        RECT 78.725 109.725 78.895 109.895 ;
        RECT 79.185 109.725 79.355 109.895 ;
        RECT 79.645 109.725 79.815 109.895 ;
        RECT 80.105 109.725 80.275 109.895 ;
        RECT 80.565 109.725 80.735 109.895 ;
        RECT 81.025 109.725 81.195 109.895 ;
        RECT 81.485 109.725 81.655 109.895 ;
        RECT 81.945 109.725 82.115 109.895 ;
        RECT 82.405 109.725 82.575 109.895 ;
        RECT 82.865 109.725 83.035 109.895 ;
        RECT 83.325 109.725 83.495 109.895 ;
        RECT 83.785 109.725 83.955 109.895 ;
        RECT 84.245 109.725 84.415 109.895 ;
        RECT 84.705 109.725 84.875 109.895 ;
        RECT 85.165 109.725 85.335 109.895 ;
        RECT 85.625 109.725 85.795 109.895 ;
        RECT 86.085 109.725 86.255 109.895 ;
        RECT 86.545 109.725 86.715 109.895 ;
        RECT 87.005 109.725 87.175 109.895 ;
        RECT 87.465 109.725 87.635 109.895 ;
        RECT 87.925 109.725 88.095 109.895 ;
        RECT 88.385 109.725 88.555 109.895 ;
        RECT 88.845 109.725 89.015 109.895 ;
        RECT 89.305 109.725 89.475 109.895 ;
        RECT 89.765 109.725 89.935 109.895 ;
        RECT 90.225 109.725 90.395 109.895 ;
        RECT 90.685 109.725 90.855 109.895 ;
        RECT 91.145 109.725 91.315 109.895 ;
        RECT 91.605 109.725 91.775 109.895 ;
        RECT 92.065 109.725 92.235 109.895 ;
        RECT 92.525 109.725 92.695 109.895 ;
        RECT 92.985 109.725 93.155 109.895 ;
        RECT 93.445 109.725 93.615 109.895 ;
        RECT 93.905 109.725 94.075 109.895 ;
        RECT 94.365 109.725 94.535 109.895 ;
        RECT 94.825 109.725 94.995 109.895 ;
        RECT 95.285 109.725 95.455 109.895 ;
        RECT 95.745 109.725 95.915 109.895 ;
        RECT 96.205 109.725 96.375 109.895 ;
        RECT 96.665 109.725 96.835 109.895 ;
        RECT 97.125 109.725 97.295 109.895 ;
        RECT 97.585 109.725 97.755 109.895 ;
        RECT 98.045 109.725 98.215 109.895 ;
        RECT 98.505 109.725 98.675 109.895 ;
        RECT 98.965 109.725 99.135 109.895 ;
        RECT 99.425 109.725 99.595 109.895 ;
        RECT 99.885 109.725 100.055 109.895 ;
        RECT 100.345 109.725 100.515 109.895 ;
        RECT 100.805 109.725 100.975 109.895 ;
        RECT 101.265 109.725 101.435 109.895 ;
        RECT 101.725 109.725 101.895 109.895 ;
        RECT 102.185 109.725 102.355 109.895 ;
        RECT 102.645 109.725 102.815 109.895 ;
        RECT 103.105 109.725 103.275 109.895 ;
        RECT 103.565 109.725 103.735 109.895 ;
        RECT 104.025 109.725 104.195 109.895 ;
        RECT 104.485 109.725 104.655 109.895 ;
        RECT 104.945 109.725 105.115 109.895 ;
        RECT 105.405 109.725 105.575 109.895 ;
        RECT 105.865 109.725 106.035 109.895 ;
        RECT 106.325 109.725 106.495 109.895 ;
        RECT 106.785 109.725 106.955 109.895 ;
        RECT 107.245 109.725 107.415 109.895 ;
        RECT 107.705 109.725 107.875 109.895 ;
        RECT 108.165 109.725 108.335 109.895 ;
        RECT 108.625 109.725 108.795 109.895 ;
        RECT 109.085 109.725 109.255 109.895 ;
        RECT 109.545 109.725 109.715 109.895 ;
        RECT 110.005 109.725 110.175 109.895 ;
        RECT 110.465 109.725 110.635 109.895 ;
        RECT 110.925 109.725 111.095 109.895 ;
        RECT 111.385 109.725 111.555 109.895 ;
        RECT 111.845 109.725 112.015 109.895 ;
        RECT 112.305 109.725 112.475 109.895 ;
        RECT 112.765 109.725 112.935 109.895 ;
        RECT 113.225 109.725 113.395 109.895 ;
        RECT 113.685 109.725 113.855 109.895 ;
        RECT 114.145 109.725 114.315 109.895 ;
        RECT 114.605 109.725 114.775 109.895 ;
        RECT 115.065 109.725 115.235 109.895 ;
        RECT 115.525 109.725 115.695 109.895 ;
        RECT 115.985 109.725 116.155 109.895 ;
        RECT 116.445 109.725 116.615 109.895 ;
        RECT 116.905 109.725 117.075 109.895 ;
        RECT 117.365 109.725 117.535 109.895 ;
        RECT 117.825 109.725 117.995 109.895 ;
        RECT 118.285 109.725 118.455 109.895 ;
        RECT 118.745 109.725 118.915 109.895 ;
        RECT 119.205 109.725 119.375 109.895 ;
        RECT 119.665 109.725 119.835 109.895 ;
        RECT 120.125 109.725 120.295 109.895 ;
        RECT 120.585 109.725 120.755 109.895 ;
        RECT 121.045 109.725 121.215 109.895 ;
        RECT 121.505 109.725 121.675 109.895 ;
        RECT 121.965 109.725 122.135 109.895 ;
        RECT 122.425 109.725 122.595 109.895 ;
        RECT 122.885 109.725 123.055 109.895 ;
        RECT 123.345 109.725 123.515 109.895 ;
        RECT 123.805 109.725 123.975 109.895 ;
        RECT 124.265 109.725 124.435 109.895 ;
        RECT 124.725 109.725 124.895 109.895 ;
        RECT 125.185 109.725 125.355 109.895 ;
        RECT 125.645 109.725 125.815 109.895 ;
        RECT 126.105 109.725 126.275 109.895 ;
        RECT 126.565 109.725 126.735 109.895 ;
        RECT 127.025 109.725 127.195 109.895 ;
        RECT 127.485 109.725 127.655 109.895 ;
        RECT 127.945 109.725 128.115 109.895 ;
        RECT 128.405 109.725 128.575 109.895 ;
        RECT 128.865 109.725 129.035 109.895 ;
        RECT 129.325 109.725 129.495 109.895 ;
        RECT 129.785 109.725 129.955 109.895 ;
        RECT 130.245 109.725 130.415 109.895 ;
        RECT 130.705 109.725 130.875 109.895 ;
        RECT 131.165 109.725 131.335 109.895 ;
        RECT 131.625 109.725 131.795 109.895 ;
        RECT 132.085 109.725 132.255 109.895 ;
        RECT 132.545 109.725 132.715 109.895 ;
        RECT 133.005 109.725 133.175 109.895 ;
        RECT 133.465 109.725 133.635 109.895 ;
        RECT 133.925 109.725 134.095 109.895 ;
        RECT 134.385 109.725 134.555 109.895 ;
        RECT 134.845 109.725 135.015 109.895 ;
        RECT 135.305 109.725 135.475 109.895 ;
        RECT 135.765 109.725 135.935 109.895 ;
        RECT 136.225 109.725 136.395 109.895 ;
        RECT 136.685 109.725 136.855 109.895 ;
        RECT 137.145 109.725 137.315 109.895 ;
        RECT 137.605 109.725 137.775 109.895 ;
        RECT 138.065 109.725 138.235 109.895 ;
        RECT 138.525 109.725 138.695 109.895 ;
        RECT 138.985 109.725 139.155 109.895 ;
        RECT 65.385 108.535 65.555 108.705 ;
        RECT 65.845 108.535 66.015 108.705 ;
        RECT 66.765 108.535 66.935 108.705 ;
        RECT 50.665 107.005 50.835 107.175 ;
        RECT 51.125 107.005 51.295 107.175 ;
        RECT 51.585 107.005 51.755 107.175 ;
        RECT 52.045 107.005 52.215 107.175 ;
        RECT 52.505 107.005 52.675 107.175 ;
        RECT 52.965 107.005 53.135 107.175 ;
        RECT 53.425 107.005 53.595 107.175 ;
        RECT 53.885 107.005 54.055 107.175 ;
        RECT 54.345 107.005 54.515 107.175 ;
        RECT 54.805 107.005 54.975 107.175 ;
        RECT 55.265 107.005 55.435 107.175 ;
        RECT 55.725 107.005 55.895 107.175 ;
        RECT 56.185 107.005 56.355 107.175 ;
        RECT 56.645 107.005 56.815 107.175 ;
        RECT 57.105 107.005 57.275 107.175 ;
        RECT 57.565 107.005 57.735 107.175 ;
        RECT 58.025 107.005 58.195 107.175 ;
        RECT 58.485 107.005 58.655 107.175 ;
        RECT 58.945 107.005 59.115 107.175 ;
        RECT 59.405 107.005 59.575 107.175 ;
        RECT 59.865 107.005 60.035 107.175 ;
        RECT 60.325 107.005 60.495 107.175 ;
        RECT 60.785 107.005 60.955 107.175 ;
        RECT 61.245 107.005 61.415 107.175 ;
        RECT 61.705 107.005 61.875 107.175 ;
        RECT 62.165 107.005 62.335 107.175 ;
        RECT 62.625 107.005 62.795 107.175 ;
        RECT 63.085 107.005 63.255 107.175 ;
        RECT 63.545 107.005 63.715 107.175 ;
        RECT 64.005 107.005 64.175 107.175 ;
        RECT 64.465 107.005 64.635 107.175 ;
        RECT 64.925 107.005 65.095 107.175 ;
        RECT 65.385 107.005 65.555 107.175 ;
        RECT 65.845 107.005 66.015 107.175 ;
        RECT 66.305 107.005 66.475 107.175 ;
        RECT 66.765 107.005 66.935 107.175 ;
        RECT 67.225 107.005 67.395 107.175 ;
        RECT 67.685 107.005 67.855 107.175 ;
        RECT 68.145 107.005 68.315 107.175 ;
        RECT 68.605 107.005 68.775 107.175 ;
        RECT 69.065 107.005 69.235 107.175 ;
        RECT 69.525 107.005 69.695 107.175 ;
        RECT 69.985 107.005 70.155 107.175 ;
        RECT 70.445 107.005 70.615 107.175 ;
        RECT 70.905 107.005 71.075 107.175 ;
        RECT 71.365 107.005 71.535 107.175 ;
        RECT 71.825 107.005 71.995 107.175 ;
        RECT 72.285 107.005 72.455 107.175 ;
        RECT 72.745 107.005 72.915 107.175 ;
        RECT 73.205 107.005 73.375 107.175 ;
        RECT 73.665 107.005 73.835 107.175 ;
        RECT 74.125 107.005 74.295 107.175 ;
        RECT 74.585 107.005 74.755 107.175 ;
        RECT 75.045 107.005 75.215 107.175 ;
        RECT 75.505 107.005 75.675 107.175 ;
        RECT 75.965 107.005 76.135 107.175 ;
        RECT 76.425 107.005 76.595 107.175 ;
        RECT 76.885 107.005 77.055 107.175 ;
        RECT 77.345 107.005 77.515 107.175 ;
        RECT 77.805 107.005 77.975 107.175 ;
        RECT 78.265 107.005 78.435 107.175 ;
        RECT 78.725 107.005 78.895 107.175 ;
        RECT 79.185 107.005 79.355 107.175 ;
        RECT 79.645 107.005 79.815 107.175 ;
        RECT 80.105 107.005 80.275 107.175 ;
        RECT 80.565 107.005 80.735 107.175 ;
        RECT 81.025 107.005 81.195 107.175 ;
        RECT 81.485 107.005 81.655 107.175 ;
        RECT 81.945 107.005 82.115 107.175 ;
        RECT 82.405 107.005 82.575 107.175 ;
        RECT 82.865 107.005 83.035 107.175 ;
        RECT 83.325 107.005 83.495 107.175 ;
        RECT 83.785 107.005 83.955 107.175 ;
        RECT 84.245 107.005 84.415 107.175 ;
        RECT 84.705 107.005 84.875 107.175 ;
        RECT 85.165 107.005 85.335 107.175 ;
        RECT 85.625 107.005 85.795 107.175 ;
        RECT 86.085 107.005 86.255 107.175 ;
        RECT 86.545 107.005 86.715 107.175 ;
        RECT 87.005 107.005 87.175 107.175 ;
        RECT 87.465 107.005 87.635 107.175 ;
        RECT 87.925 107.005 88.095 107.175 ;
        RECT 88.385 107.005 88.555 107.175 ;
        RECT 88.845 107.005 89.015 107.175 ;
        RECT 89.305 107.005 89.475 107.175 ;
        RECT 89.765 107.005 89.935 107.175 ;
        RECT 90.225 107.005 90.395 107.175 ;
        RECT 90.685 107.005 90.855 107.175 ;
        RECT 91.145 107.005 91.315 107.175 ;
        RECT 91.605 107.005 91.775 107.175 ;
        RECT 92.065 107.005 92.235 107.175 ;
        RECT 92.525 107.005 92.695 107.175 ;
        RECT 92.985 107.005 93.155 107.175 ;
        RECT 93.445 107.005 93.615 107.175 ;
        RECT 93.905 107.005 94.075 107.175 ;
        RECT 94.365 107.005 94.535 107.175 ;
        RECT 94.825 107.005 94.995 107.175 ;
        RECT 95.285 107.005 95.455 107.175 ;
        RECT 95.745 107.005 95.915 107.175 ;
        RECT 96.205 107.005 96.375 107.175 ;
        RECT 96.665 107.005 96.835 107.175 ;
        RECT 97.125 107.005 97.295 107.175 ;
        RECT 97.585 107.005 97.755 107.175 ;
        RECT 98.045 107.005 98.215 107.175 ;
        RECT 98.505 107.005 98.675 107.175 ;
        RECT 98.965 107.005 99.135 107.175 ;
        RECT 99.425 107.005 99.595 107.175 ;
        RECT 99.885 107.005 100.055 107.175 ;
        RECT 100.345 107.005 100.515 107.175 ;
        RECT 100.805 107.005 100.975 107.175 ;
        RECT 101.265 107.005 101.435 107.175 ;
        RECT 101.725 107.005 101.895 107.175 ;
        RECT 102.185 107.005 102.355 107.175 ;
        RECT 102.645 107.005 102.815 107.175 ;
        RECT 103.105 107.005 103.275 107.175 ;
        RECT 103.565 107.005 103.735 107.175 ;
        RECT 104.025 107.005 104.195 107.175 ;
        RECT 104.485 107.005 104.655 107.175 ;
        RECT 104.945 107.005 105.115 107.175 ;
        RECT 105.405 107.005 105.575 107.175 ;
        RECT 105.865 107.005 106.035 107.175 ;
        RECT 106.325 107.005 106.495 107.175 ;
        RECT 106.785 107.005 106.955 107.175 ;
        RECT 107.245 107.005 107.415 107.175 ;
        RECT 107.705 107.005 107.875 107.175 ;
        RECT 108.165 107.005 108.335 107.175 ;
        RECT 108.625 107.005 108.795 107.175 ;
        RECT 109.085 107.005 109.255 107.175 ;
        RECT 109.545 107.005 109.715 107.175 ;
        RECT 110.005 107.005 110.175 107.175 ;
        RECT 110.465 107.005 110.635 107.175 ;
        RECT 110.925 107.005 111.095 107.175 ;
        RECT 111.385 107.005 111.555 107.175 ;
        RECT 111.845 107.005 112.015 107.175 ;
        RECT 112.305 107.005 112.475 107.175 ;
        RECT 112.765 107.005 112.935 107.175 ;
        RECT 113.225 107.005 113.395 107.175 ;
        RECT 113.685 107.005 113.855 107.175 ;
        RECT 114.145 107.005 114.315 107.175 ;
        RECT 114.605 107.005 114.775 107.175 ;
        RECT 115.065 107.005 115.235 107.175 ;
        RECT 115.525 107.005 115.695 107.175 ;
        RECT 115.985 107.005 116.155 107.175 ;
        RECT 116.445 107.005 116.615 107.175 ;
        RECT 116.905 107.005 117.075 107.175 ;
        RECT 117.365 107.005 117.535 107.175 ;
        RECT 117.825 107.005 117.995 107.175 ;
        RECT 118.285 107.005 118.455 107.175 ;
        RECT 118.745 107.005 118.915 107.175 ;
        RECT 119.205 107.005 119.375 107.175 ;
        RECT 119.665 107.005 119.835 107.175 ;
        RECT 120.125 107.005 120.295 107.175 ;
        RECT 120.585 107.005 120.755 107.175 ;
        RECT 121.045 107.005 121.215 107.175 ;
        RECT 121.505 107.005 121.675 107.175 ;
        RECT 121.965 107.005 122.135 107.175 ;
        RECT 122.425 107.005 122.595 107.175 ;
        RECT 122.885 107.005 123.055 107.175 ;
        RECT 123.345 107.005 123.515 107.175 ;
        RECT 123.805 107.005 123.975 107.175 ;
        RECT 124.265 107.005 124.435 107.175 ;
        RECT 124.725 107.005 124.895 107.175 ;
        RECT 125.185 107.005 125.355 107.175 ;
        RECT 125.645 107.005 125.815 107.175 ;
        RECT 126.105 107.005 126.275 107.175 ;
        RECT 126.565 107.005 126.735 107.175 ;
        RECT 127.025 107.005 127.195 107.175 ;
        RECT 127.485 107.005 127.655 107.175 ;
        RECT 127.945 107.005 128.115 107.175 ;
        RECT 128.405 107.005 128.575 107.175 ;
        RECT 128.865 107.005 129.035 107.175 ;
        RECT 129.325 107.005 129.495 107.175 ;
        RECT 129.785 107.005 129.955 107.175 ;
        RECT 130.245 107.005 130.415 107.175 ;
        RECT 130.705 107.005 130.875 107.175 ;
        RECT 131.165 107.005 131.335 107.175 ;
        RECT 131.625 107.005 131.795 107.175 ;
        RECT 132.085 107.005 132.255 107.175 ;
        RECT 132.545 107.005 132.715 107.175 ;
        RECT 133.005 107.005 133.175 107.175 ;
        RECT 133.465 107.005 133.635 107.175 ;
        RECT 133.925 107.005 134.095 107.175 ;
        RECT 134.385 107.005 134.555 107.175 ;
        RECT 134.845 107.005 135.015 107.175 ;
        RECT 135.305 107.005 135.475 107.175 ;
        RECT 135.765 107.005 135.935 107.175 ;
        RECT 136.225 107.005 136.395 107.175 ;
        RECT 136.685 107.005 136.855 107.175 ;
        RECT 137.145 107.005 137.315 107.175 ;
        RECT 137.605 107.005 137.775 107.175 ;
        RECT 138.065 107.005 138.235 107.175 ;
        RECT 138.525 107.005 138.695 107.175 ;
        RECT 138.985 107.005 139.155 107.175 ;
        RECT 58.025 105.815 58.195 105.985 ;
        RECT 57.105 105.475 57.275 105.645 ;
        RECT 57.565 105.475 57.735 105.645 ;
        RECT 58.485 105.475 58.655 105.645 ;
        RECT 61.245 105.815 61.415 105.985 ;
        RECT 58.945 105.135 59.115 105.305 ;
        RECT 62.165 105.475 62.335 105.645 ;
        RECT 50.665 104.285 50.835 104.455 ;
        RECT 51.125 104.285 51.295 104.455 ;
        RECT 51.585 104.285 51.755 104.455 ;
        RECT 52.045 104.285 52.215 104.455 ;
        RECT 52.505 104.285 52.675 104.455 ;
        RECT 52.965 104.285 53.135 104.455 ;
        RECT 53.425 104.285 53.595 104.455 ;
        RECT 53.885 104.285 54.055 104.455 ;
        RECT 54.345 104.285 54.515 104.455 ;
        RECT 54.805 104.285 54.975 104.455 ;
        RECT 55.265 104.285 55.435 104.455 ;
        RECT 55.725 104.285 55.895 104.455 ;
        RECT 56.185 104.285 56.355 104.455 ;
        RECT 56.645 104.285 56.815 104.455 ;
        RECT 57.105 104.285 57.275 104.455 ;
        RECT 57.565 104.285 57.735 104.455 ;
        RECT 58.025 104.285 58.195 104.455 ;
        RECT 58.485 104.285 58.655 104.455 ;
        RECT 58.945 104.285 59.115 104.455 ;
        RECT 59.405 104.285 59.575 104.455 ;
        RECT 59.865 104.285 60.035 104.455 ;
        RECT 60.325 104.285 60.495 104.455 ;
        RECT 60.785 104.285 60.955 104.455 ;
        RECT 61.245 104.285 61.415 104.455 ;
        RECT 61.705 104.285 61.875 104.455 ;
        RECT 62.165 104.285 62.335 104.455 ;
        RECT 62.625 104.285 62.795 104.455 ;
        RECT 63.085 104.285 63.255 104.455 ;
        RECT 63.545 104.285 63.715 104.455 ;
        RECT 64.005 104.285 64.175 104.455 ;
        RECT 64.465 104.285 64.635 104.455 ;
        RECT 64.925 104.285 65.095 104.455 ;
        RECT 65.385 104.285 65.555 104.455 ;
        RECT 65.845 104.285 66.015 104.455 ;
        RECT 66.305 104.285 66.475 104.455 ;
        RECT 66.765 104.285 66.935 104.455 ;
        RECT 67.225 104.285 67.395 104.455 ;
        RECT 67.685 104.285 67.855 104.455 ;
        RECT 68.145 104.285 68.315 104.455 ;
        RECT 68.605 104.285 68.775 104.455 ;
        RECT 69.065 104.285 69.235 104.455 ;
        RECT 69.525 104.285 69.695 104.455 ;
        RECT 69.985 104.285 70.155 104.455 ;
        RECT 70.445 104.285 70.615 104.455 ;
        RECT 70.905 104.285 71.075 104.455 ;
        RECT 71.365 104.285 71.535 104.455 ;
        RECT 71.825 104.285 71.995 104.455 ;
        RECT 72.285 104.285 72.455 104.455 ;
        RECT 72.745 104.285 72.915 104.455 ;
        RECT 73.205 104.285 73.375 104.455 ;
        RECT 73.665 104.285 73.835 104.455 ;
        RECT 74.125 104.285 74.295 104.455 ;
        RECT 74.585 104.285 74.755 104.455 ;
        RECT 75.045 104.285 75.215 104.455 ;
        RECT 75.505 104.285 75.675 104.455 ;
        RECT 75.965 104.285 76.135 104.455 ;
        RECT 76.425 104.285 76.595 104.455 ;
        RECT 76.885 104.285 77.055 104.455 ;
        RECT 77.345 104.285 77.515 104.455 ;
        RECT 77.805 104.285 77.975 104.455 ;
        RECT 78.265 104.285 78.435 104.455 ;
        RECT 78.725 104.285 78.895 104.455 ;
        RECT 79.185 104.285 79.355 104.455 ;
        RECT 79.645 104.285 79.815 104.455 ;
        RECT 80.105 104.285 80.275 104.455 ;
        RECT 80.565 104.285 80.735 104.455 ;
        RECT 81.025 104.285 81.195 104.455 ;
        RECT 81.485 104.285 81.655 104.455 ;
        RECT 81.945 104.285 82.115 104.455 ;
        RECT 82.405 104.285 82.575 104.455 ;
        RECT 82.865 104.285 83.035 104.455 ;
        RECT 83.325 104.285 83.495 104.455 ;
        RECT 83.785 104.285 83.955 104.455 ;
        RECT 84.245 104.285 84.415 104.455 ;
        RECT 84.705 104.285 84.875 104.455 ;
        RECT 85.165 104.285 85.335 104.455 ;
        RECT 85.625 104.285 85.795 104.455 ;
        RECT 86.085 104.285 86.255 104.455 ;
        RECT 86.545 104.285 86.715 104.455 ;
        RECT 87.005 104.285 87.175 104.455 ;
        RECT 87.465 104.285 87.635 104.455 ;
        RECT 87.925 104.285 88.095 104.455 ;
        RECT 88.385 104.285 88.555 104.455 ;
        RECT 88.845 104.285 89.015 104.455 ;
        RECT 89.305 104.285 89.475 104.455 ;
        RECT 89.765 104.285 89.935 104.455 ;
        RECT 90.225 104.285 90.395 104.455 ;
        RECT 90.685 104.285 90.855 104.455 ;
        RECT 91.145 104.285 91.315 104.455 ;
        RECT 91.605 104.285 91.775 104.455 ;
        RECT 92.065 104.285 92.235 104.455 ;
        RECT 92.525 104.285 92.695 104.455 ;
        RECT 92.985 104.285 93.155 104.455 ;
        RECT 93.445 104.285 93.615 104.455 ;
        RECT 93.905 104.285 94.075 104.455 ;
        RECT 94.365 104.285 94.535 104.455 ;
        RECT 94.825 104.285 94.995 104.455 ;
        RECT 95.285 104.285 95.455 104.455 ;
        RECT 95.745 104.285 95.915 104.455 ;
        RECT 96.205 104.285 96.375 104.455 ;
        RECT 96.665 104.285 96.835 104.455 ;
        RECT 97.125 104.285 97.295 104.455 ;
        RECT 97.585 104.285 97.755 104.455 ;
        RECT 98.045 104.285 98.215 104.455 ;
        RECT 98.505 104.285 98.675 104.455 ;
        RECT 98.965 104.285 99.135 104.455 ;
        RECT 99.425 104.285 99.595 104.455 ;
        RECT 99.885 104.285 100.055 104.455 ;
        RECT 100.345 104.285 100.515 104.455 ;
        RECT 100.805 104.285 100.975 104.455 ;
        RECT 101.265 104.285 101.435 104.455 ;
        RECT 101.725 104.285 101.895 104.455 ;
        RECT 102.185 104.285 102.355 104.455 ;
        RECT 102.645 104.285 102.815 104.455 ;
        RECT 103.105 104.285 103.275 104.455 ;
        RECT 103.565 104.285 103.735 104.455 ;
        RECT 104.025 104.285 104.195 104.455 ;
        RECT 104.485 104.285 104.655 104.455 ;
        RECT 104.945 104.285 105.115 104.455 ;
        RECT 105.405 104.285 105.575 104.455 ;
        RECT 105.865 104.285 106.035 104.455 ;
        RECT 106.325 104.285 106.495 104.455 ;
        RECT 106.785 104.285 106.955 104.455 ;
        RECT 107.245 104.285 107.415 104.455 ;
        RECT 107.705 104.285 107.875 104.455 ;
        RECT 108.165 104.285 108.335 104.455 ;
        RECT 108.625 104.285 108.795 104.455 ;
        RECT 109.085 104.285 109.255 104.455 ;
        RECT 109.545 104.285 109.715 104.455 ;
        RECT 110.005 104.285 110.175 104.455 ;
        RECT 110.465 104.285 110.635 104.455 ;
        RECT 110.925 104.285 111.095 104.455 ;
        RECT 111.385 104.285 111.555 104.455 ;
        RECT 111.845 104.285 112.015 104.455 ;
        RECT 112.305 104.285 112.475 104.455 ;
        RECT 112.765 104.285 112.935 104.455 ;
        RECT 113.225 104.285 113.395 104.455 ;
        RECT 113.685 104.285 113.855 104.455 ;
        RECT 114.145 104.285 114.315 104.455 ;
        RECT 114.605 104.285 114.775 104.455 ;
        RECT 115.065 104.285 115.235 104.455 ;
        RECT 115.525 104.285 115.695 104.455 ;
        RECT 115.985 104.285 116.155 104.455 ;
        RECT 116.445 104.285 116.615 104.455 ;
        RECT 116.905 104.285 117.075 104.455 ;
        RECT 117.365 104.285 117.535 104.455 ;
        RECT 117.825 104.285 117.995 104.455 ;
        RECT 118.285 104.285 118.455 104.455 ;
        RECT 118.745 104.285 118.915 104.455 ;
        RECT 119.205 104.285 119.375 104.455 ;
        RECT 119.665 104.285 119.835 104.455 ;
        RECT 120.125 104.285 120.295 104.455 ;
        RECT 120.585 104.285 120.755 104.455 ;
        RECT 121.045 104.285 121.215 104.455 ;
        RECT 121.505 104.285 121.675 104.455 ;
        RECT 121.965 104.285 122.135 104.455 ;
        RECT 122.425 104.285 122.595 104.455 ;
        RECT 122.885 104.285 123.055 104.455 ;
        RECT 123.345 104.285 123.515 104.455 ;
        RECT 123.805 104.285 123.975 104.455 ;
        RECT 124.265 104.285 124.435 104.455 ;
        RECT 124.725 104.285 124.895 104.455 ;
        RECT 125.185 104.285 125.355 104.455 ;
        RECT 125.645 104.285 125.815 104.455 ;
        RECT 126.105 104.285 126.275 104.455 ;
        RECT 126.565 104.285 126.735 104.455 ;
        RECT 127.025 104.285 127.195 104.455 ;
        RECT 127.485 104.285 127.655 104.455 ;
        RECT 127.945 104.285 128.115 104.455 ;
        RECT 128.405 104.285 128.575 104.455 ;
        RECT 128.865 104.285 129.035 104.455 ;
        RECT 129.325 104.285 129.495 104.455 ;
        RECT 129.785 104.285 129.955 104.455 ;
        RECT 130.245 104.285 130.415 104.455 ;
        RECT 130.705 104.285 130.875 104.455 ;
        RECT 131.165 104.285 131.335 104.455 ;
        RECT 131.625 104.285 131.795 104.455 ;
        RECT 132.085 104.285 132.255 104.455 ;
        RECT 132.545 104.285 132.715 104.455 ;
        RECT 133.005 104.285 133.175 104.455 ;
        RECT 133.465 104.285 133.635 104.455 ;
        RECT 133.925 104.285 134.095 104.455 ;
        RECT 134.385 104.285 134.555 104.455 ;
        RECT 134.845 104.285 135.015 104.455 ;
        RECT 135.305 104.285 135.475 104.455 ;
        RECT 135.765 104.285 135.935 104.455 ;
        RECT 136.225 104.285 136.395 104.455 ;
        RECT 136.685 104.285 136.855 104.455 ;
        RECT 137.145 104.285 137.315 104.455 ;
        RECT 137.605 104.285 137.775 104.455 ;
        RECT 138.065 104.285 138.235 104.455 ;
        RECT 138.525 104.285 138.695 104.455 ;
        RECT 138.985 104.285 139.155 104.455 ;
        RECT 52.965 103.775 53.135 103.945 ;
        RECT 52.045 103.095 52.215 103.265 ;
        RECT 61.705 103.435 61.875 103.605 ;
        RECT 59.865 103.095 60.035 103.265 ;
        RECT 61.245 103.095 61.415 103.265 ;
        RECT 62.170 103.095 62.340 103.265 ;
        RECT 63.085 103.435 63.255 103.605 ;
        RECT 65.400 103.095 65.570 103.265 ;
        RECT 62.625 102.755 62.795 102.925 ;
        RECT 64.005 102.755 64.175 102.925 ;
        RECT 50.665 101.565 50.835 101.735 ;
        RECT 51.125 101.565 51.295 101.735 ;
        RECT 51.585 101.565 51.755 101.735 ;
        RECT 52.045 101.565 52.215 101.735 ;
        RECT 52.505 101.565 52.675 101.735 ;
        RECT 52.965 101.565 53.135 101.735 ;
        RECT 53.425 101.565 53.595 101.735 ;
        RECT 53.885 101.565 54.055 101.735 ;
        RECT 54.345 101.565 54.515 101.735 ;
        RECT 54.805 101.565 54.975 101.735 ;
        RECT 55.265 101.565 55.435 101.735 ;
        RECT 55.725 101.565 55.895 101.735 ;
        RECT 56.185 101.565 56.355 101.735 ;
        RECT 56.645 101.565 56.815 101.735 ;
        RECT 57.105 101.565 57.275 101.735 ;
        RECT 57.565 101.565 57.735 101.735 ;
        RECT 58.025 101.565 58.195 101.735 ;
        RECT 58.485 101.565 58.655 101.735 ;
        RECT 58.945 101.565 59.115 101.735 ;
        RECT 59.405 101.565 59.575 101.735 ;
        RECT 59.865 101.565 60.035 101.735 ;
        RECT 60.325 101.565 60.495 101.735 ;
        RECT 60.785 101.565 60.955 101.735 ;
        RECT 61.245 101.565 61.415 101.735 ;
        RECT 61.705 101.565 61.875 101.735 ;
        RECT 62.165 101.565 62.335 101.735 ;
        RECT 62.625 101.565 62.795 101.735 ;
        RECT 63.085 101.565 63.255 101.735 ;
        RECT 63.545 101.565 63.715 101.735 ;
        RECT 64.005 101.565 64.175 101.735 ;
        RECT 64.465 101.565 64.635 101.735 ;
        RECT 64.925 101.565 65.095 101.735 ;
        RECT 65.385 101.565 65.555 101.735 ;
        RECT 65.845 101.565 66.015 101.735 ;
        RECT 66.305 101.565 66.475 101.735 ;
        RECT 66.765 101.565 66.935 101.735 ;
        RECT 67.225 101.565 67.395 101.735 ;
        RECT 67.685 101.565 67.855 101.735 ;
        RECT 68.145 101.565 68.315 101.735 ;
        RECT 68.605 101.565 68.775 101.735 ;
        RECT 69.065 101.565 69.235 101.735 ;
        RECT 69.525 101.565 69.695 101.735 ;
        RECT 69.985 101.565 70.155 101.735 ;
        RECT 70.445 101.565 70.615 101.735 ;
        RECT 70.905 101.565 71.075 101.735 ;
        RECT 71.365 101.565 71.535 101.735 ;
        RECT 71.825 101.565 71.995 101.735 ;
        RECT 72.285 101.565 72.455 101.735 ;
        RECT 72.745 101.565 72.915 101.735 ;
        RECT 73.205 101.565 73.375 101.735 ;
        RECT 73.665 101.565 73.835 101.735 ;
        RECT 74.125 101.565 74.295 101.735 ;
        RECT 74.585 101.565 74.755 101.735 ;
        RECT 75.045 101.565 75.215 101.735 ;
        RECT 75.505 101.565 75.675 101.735 ;
        RECT 75.965 101.565 76.135 101.735 ;
        RECT 76.425 101.565 76.595 101.735 ;
        RECT 76.885 101.565 77.055 101.735 ;
        RECT 77.345 101.565 77.515 101.735 ;
        RECT 77.805 101.565 77.975 101.735 ;
        RECT 78.265 101.565 78.435 101.735 ;
        RECT 78.725 101.565 78.895 101.735 ;
        RECT 79.185 101.565 79.355 101.735 ;
        RECT 79.645 101.565 79.815 101.735 ;
        RECT 80.105 101.565 80.275 101.735 ;
        RECT 80.565 101.565 80.735 101.735 ;
        RECT 81.025 101.565 81.195 101.735 ;
        RECT 81.485 101.565 81.655 101.735 ;
        RECT 81.945 101.565 82.115 101.735 ;
        RECT 82.405 101.565 82.575 101.735 ;
        RECT 82.865 101.565 83.035 101.735 ;
        RECT 83.325 101.565 83.495 101.735 ;
        RECT 83.785 101.565 83.955 101.735 ;
        RECT 84.245 101.565 84.415 101.735 ;
        RECT 84.705 101.565 84.875 101.735 ;
        RECT 85.165 101.565 85.335 101.735 ;
        RECT 85.625 101.565 85.795 101.735 ;
        RECT 86.085 101.565 86.255 101.735 ;
        RECT 86.545 101.565 86.715 101.735 ;
        RECT 87.005 101.565 87.175 101.735 ;
        RECT 87.465 101.565 87.635 101.735 ;
        RECT 87.925 101.565 88.095 101.735 ;
        RECT 88.385 101.565 88.555 101.735 ;
        RECT 88.845 101.565 89.015 101.735 ;
        RECT 89.305 101.565 89.475 101.735 ;
        RECT 89.765 101.565 89.935 101.735 ;
        RECT 90.225 101.565 90.395 101.735 ;
        RECT 90.685 101.565 90.855 101.735 ;
        RECT 91.145 101.565 91.315 101.735 ;
        RECT 91.605 101.565 91.775 101.735 ;
        RECT 92.065 101.565 92.235 101.735 ;
        RECT 92.525 101.565 92.695 101.735 ;
        RECT 92.985 101.565 93.155 101.735 ;
        RECT 93.445 101.565 93.615 101.735 ;
        RECT 93.905 101.565 94.075 101.735 ;
        RECT 94.365 101.565 94.535 101.735 ;
        RECT 94.825 101.565 94.995 101.735 ;
        RECT 95.285 101.565 95.455 101.735 ;
        RECT 95.745 101.565 95.915 101.735 ;
        RECT 96.205 101.565 96.375 101.735 ;
        RECT 96.665 101.565 96.835 101.735 ;
        RECT 97.125 101.565 97.295 101.735 ;
        RECT 97.585 101.565 97.755 101.735 ;
        RECT 98.045 101.565 98.215 101.735 ;
        RECT 98.505 101.565 98.675 101.735 ;
        RECT 98.965 101.565 99.135 101.735 ;
        RECT 99.425 101.565 99.595 101.735 ;
        RECT 99.885 101.565 100.055 101.735 ;
        RECT 100.345 101.565 100.515 101.735 ;
        RECT 100.805 101.565 100.975 101.735 ;
        RECT 101.265 101.565 101.435 101.735 ;
        RECT 101.725 101.565 101.895 101.735 ;
        RECT 102.185 101.565 102.355 101.735 ;
        RECT 102.645 101.565 102.815 101.735 ;
        RECT 103.105 101.565 103.275 101.735 ;
        RECT 103.565 101.565 103.735 101.735 ;
        RECT 104.025 101.565 104.195 101.735 ;
        RECT 104.485 101.565 104.655 101.735 ;
        RECT 104.945 101.565 105.115 101.735 ;
        RECT 105.405 101.565 105.575 101.735 ;
        RECT 105.865 101.565 106.035 101.735 ;
        RECT 106.325 101.565 106.495 101.735 ;
        RECT 106.785 101.565 106.955 101.735 ;
        RECT 107.245 101.565 107.415 101.735 ;
        RECT 107.705 101.565 107.875 101.735 ;
        RECT 108.165 101.565 108.335 101.735 ;
        RECT 108.625 101.565 108.795 101.735 ;
        RECT 109.085 101.565 109.255 101.735 ;
        RECT 109.545 101.565 109.715 101.735 ;
        RECT 110.005 101.565 110.175 101.735 ;
        RECT 110.465 101.565 110.635 101.735 ;
        RECT 110.925 101.565 111.095 101.735 ;
        RECT 111.385 101.565 111.555 101.735 ;
        RECT 111.845 101.565 112.015 101.735 ;
        RECT 112.305 101.565 112.475 101.735 ;
        RECT 112.765 101.565 112.935 101.735 ;
        RECT 113.225 101.565 113.395 101.735 ;
        RECT 113.685 101.565 113.855 101.735 ;
        RECT 114.145 101.565 114.315 101.735 ;
        RECT 114.605 101.565 114.775 101.735 ;
        RECT 115.065 101.565 115.235 101.735 ;
        RECT 115.525 101.565 115.695 101.735 ;
        RECT 115.985 101.565 116.155 101.735 ;
        RECT 116.445 101.565 116.615 101.735 ;
        RECT 116.905 101.565 117.075 101.735 ;
        RECT 117.365 101.565 117.535 101.735 ;
        RECT 117.825 101.565 117.995 101.735 ;
        RECT 118.285 101.565 118.455 101.735 ;
        RECT 118.745 101.565 118.915 101.735 ;
        RECT 119.205 101.565 119.375 101.735 ;
        RECT 119.665 101.565 119.835 101.735 ;
        RECT 120.125 101.565 120.295 101.735 ;
        RECT 120.585 101.565 120.755 101.735 ;
        RECT 121.045 101.565 121.215 101.735 ;
        RECT 121.505 101.565 121.675 101.735 ;
        RECT 121.965 101.565 122.135 101.735 ;
        RECT 122.425 101.565 122.595 101.735 ;
        RECT 122.885 101.565 123.055 101.735 ;
        RECT 123.345 101.565 123.515 101.735 ;
        RECT 123.805 101.565 123.975 101.735 ;
        RECT 124.265 101.565 124.435 101.735 ;
        RECT 124.725 101.565 124.895 101.735 ;
        RECT 125.185 101.565 125.355 101.735 ;
        RECT 125.645 101.565 125.815 101.735 ;
        RECT 126.105 101.565 126.275 101.735 ;
        RECT 126.565 101.565 126.735 101.735 ;
        RECT 127.025 101.565 127.195 101.735 ;
        RECT 127.485 101.565 127.655 101.735 ;
        RECT 127.945 101.565 128.115 101.735 ;
        RECT 128.405 101.565 128.575 101.735 ;
        RECT 128.865 101.565 129.035 101.735 ;
        RECT 129.325 101.565 129.495 101.735 ;
        RECT 129.785 101.565 129.955 101.735 ;
        RECT 130.245 101.565 130.415 101.735 ;
        RECT 130.705 101.565 130.875 101.735 ;
        RECT 131.165 101.565 131.335 101.735 ;
        RECT 131.625 101.565 131.795 101.735 ;
        RECT 132.085 101.565 132.255 101.735 ;
        RECT 132.545 101.565 132.715 101.735 ;
        RECT 133.005 101.565 133.175 101.735 ;
        RECT 133.465 101.565 133.635 101.735 ;
        RECT 133.925 101.565 134.095 101.735 ;
        RECT 134.385 101.565 134.555 101.735 ;
        RECT 134.845 101.565 135.015 101.735 ;
        RECT 135.305 101.565 135.475 101.735 ;
        RECT 135.765 101.565 135.935 101.735 ;
        RECT 136.225 101.565 136.395 101.735 ;
        RECT 136.685 101.565 136.855 101.735 ;
        RECT 137.145 101.565 137.315 101.735 ;
        RECT 137.605 101.565 137.775 101.735 ;
        RECT 138.065 101.565 138.235 101.735 ;
        RECT 138.525 101.565 138.695 101.735 ;
        RECT 138.985 101.565 139.155 101.735 ;
        RECT 52.045 100.035 52.215 100.205 ;
        RECT 52.965 99.355 53.135 99.525 ;
        RECT 50.665 98.845 50.835 99.015 ;
        RECT 51.125 98.845 51.295 99.015 ;
        RECT 51.585 98.845 51.755 99.015 ;
        RECT 52.045 98.845 52.215 99.015 ;
        RECT 52.505 98.845 52.675 99.015 ;
        RECT 52.965 98.845 53.135 99.015 ;
        RECT 53.425 98.845 53.595 99.015 ;
        RECT 53.885 98.845 54.055 99.015 ;
        RECT 54.345 98.845 54.515 99.015 ;
        RECT 54.805 98.845 54.975 99.015 ;
        RECT 55.265 98.845 55.435 99.015 ;
        RECT 55.725 98.845 55.895 99.015 ;
        RECT 56.185 98.845 56.355 99.015 ;
        RECT 56.645 98.845 56.815 99.015 ;
        RECT 57.105 98.845 57.275 99.015 ;
        RECT 57.565 98.845 57.735 99.015 ;
        RECT 58.025 98.845 58.195 99.015 ;
        RECT 58.485 98.845 58.655 99.015 ;
        RECT 58.945 98.845 59.115 99.015 ;
        RECT 59.405 98.845 59.575 99.015 ;
        RECT 59.865 98.845 60.035 99.015 ;
        RECT 60.325 98.845 60.495 99.015 ;
        RECT 60.785 98.845 60.955 99.015 ;
        RECT 61.245 98.845 61.415 99.015 ;
        RECT 61.705 98.845 61.875 99.015 ;
        RECT 62.165 98.845 62.335 99.015 ;
        RECT 62.625 98.845 62.795 99.015 ;
        RECT 63.085 98.845 63.255 99.015 ;
        RECT 63.545 98.845 63.715 99.015 ;
        RECT 64.005 98.845 64.175 99.015 ;
        RECT 64.465 98.845 64.635 99.015 ;
        RECT 64.925 98.845 65.095 99.015 ;
        RECT 65.385 98.845 65.555 99.015 ;
        RECT 65.845 98.845 66.015 99.015 ;
        RECT 66.305 98.845 66.475 99.015 ;
        RECT 66.765 98.845 66.935 99.015 ;
        RECT 67.225 98.845 67.395 99.015 ;
        RECT 67.685 98.845 67.855 99.015 ;
        RECT 68.145 98.845 68.315 99.015 ;
        RECT 68.605 98.845 68.775 99.015 ;
        RECT 69.065 98.845 69.235 99.015 ;
        RECT 69.525 98.845 69.695 99.015 ;
        RECT 69.985 98.845 70.155 99.015 ;
        RECT 70.445 98.845 70.615 99.015 ;
        RECT 70.905 98.845 71.075 99.015 ;
        RECT 71.365 98.845 71.535 99.015 ;
        RECT 71.825 98.845 71.995 99.015 ;
        RECT 72.285 98.845 72.455 99.015 ;
        RECT 72.745 98.845 72.915 99.015 ;
        RECT 73.205 98.845 73.375 99.015 ;
        RECT 73.665 98.845 73.835 99.015 ;
        RECT 74.125 98.845 74.295 99.015 ;
        RECT 74.585 98.845 74.755 99.015 ;
        RECT 75.045 98.845 75.215 99.015 ;
        RECT 75.505 98.845 75.675 99.015 ;
        RECT 75.965 98.845 76.135 99.015 ;
        RECT 76.425 98.845 76.595 99.015 ;
        RECT 76.885 98.845 77.055 99.015 ;
        RECT 77.345 98.845 77.515 99.015 ;
        RECT 77.805 98.845 77.975 99.015 ;
        RECT 78.265 98.845 78.435 99.015 ;
        RECT 78.725 98.845 78.895 99.015 ;
        RECT 79.185 98.845 79.355 99.015 ;
        RECT 79.645 98.845 79.815 99.015 ;
        RECT 80.105 98.845 80.275 99.015 ;
        RECT 80.565 98.845 80.735 99.015 ;
        RECT 81.025 98.845 81.195 99.015 ;
        RECT 81.485 98.845 81.655 99.015 ;
        RECT 81.945 98.845 82.115 99.015 ;
        RECT 82.405 98.845 82.575 99.015 ;
        RECT 82.865 98.845 83.035 99.015 ;
        RECT 83.325 98.845 83.495 99.015 ;
        RECT 83.785 98.845 83.955 99.015 ;
        RECT 84.245 98.845 84.415 99.015 ;
        RECT 84.705 98.845 84.875 99.015 ;
        RECT 85.165 98.845 85.335 99.015 ;
        RECT 85.625 98.845 85.795 99.015 ;
        RECT 86.085 98.845 86.255 99.015 ;
        RECT 86.545 98.845 86.715 99.015 ;
        RECT 87.005 98.845 87.175 99.015 ;
        RECT 87.465 98.845 87.635 99.015 ;
        RECT 87.925 98.845 88.095 99.015 ;
        RECT 88.385 98.845 88.555 99.015 ;
        RECT 88.845 98.845 89.015 99.015 ;
        RECT 89.305 98.845 89.475 99.015 ;
        RECT 89.765 98.845 89.935 99.015 ;
        RECT 90.225 98.845 90.395 99.015 ;
        RECT 90.685 98.845 90.855 99.015 ;
        RECT 91.145 98.845 91.315 99.015 ;
        RECT 91.605 98.845 91.775 99.015 ;
        RECT 92.065 98.845 92.235 99.015 ;
        RECT 92.525 98.845 92.695 99.015 ;
        RECT 92.985 98.845 93.155 99.015 ;
        RECT 93.445 98.845 93.615 99.015 ;
        RECT 93.905 98.845 94.075 99.015 ;
        RECT 94.365 98.845 94.535 99.015 ;
        RECT 94.825 98.845 94.995 99.015 ;
        RECT 95.285 98.845 95.455 99.015 ;
        RECT 95.745 98.845 95.915 99.015 ;
        RECT 96.205 98.845 96.375 99.015 ;
        RECT 96.665 98.845 96.835 99.015 ;
        RECT 97.125 98.845 97.295 99.015 ;
        RECT 97.585 98.845 97.755 99.015 ;
        RECT 98.045 98.845 98.215 99.015 ;
        RECT 98.505 98.845 98.675 99.015 ;
        RECT 98.965 98.845 99.135 99.015 ;
        RECT 99.425 98.845 99.595 99.015 ;
        RECT 99.885 98.845 100.055 99.015 ;
        RECT 100.345 98.845 100.515 99.015 ;
        RECT 100.805 98.845 100.975 99.015 ;
        RECT 101.265 98.845 101.435 99.015 ;
        RECT 101.725 98.845 101.895 99.015 ;
        RECT 102.185 98.845 102.355 99.015 ;
        RECT 102.645 98.845 102.815 99.015 ;
        RECT 103.105 98.845 103.275 99.015 ;
        RECT 103.565 98.845 103.735 99.015 ;
        RECT 104.025 98.845 104.195 99.015 ;
        RECT 104.485 98.845 104.655 99.015 ;
        RECT 104.945 98.845 105.115 99.015 ;
        RECT 105.405 98.845 105.575 99.015 ;
        RECT 105.865 98.845 106.035 99.015 ;
        RECT 106.325 98.845 106.495 99.015 ;
        RECT 106.785 98.845 106.955 99.015 ;
        RECT 107.245 98.845 107.415 99.015 ;
        RECT 107.705 98.845 107.875 99.015 ;
        RECT 108.165 98.845 108.335 99.015 ;
        RECT 108.625 98.845 108.795 99.015 ;
        RECT 109.085 98.845 109.255 99.015 ;
        RECT 109.545 98.845 109.715 99.015 ;
        RECT 110.005 98.845 110.175 99.015 ;
        RECT 110.465 98.845 110.635 99.015 ;
        RECT 110.925 98.845 111.095 99.015 ;
        RECT 111.385 98.845 111.555 99.015 ;
        RECT 111.845 98.845 112.015 99.015 ;
        RECT 112.305 98.845 112.475 99.015 ;
        RECT 112.765 98.845 112.935 99.015 ;
        RECT 113.225 98.845 113.395 99.015 ;
        RECT 113.685 98.845 113.855 99.015 ;
        RECT 114.145 98.845 114.315 99.015 ;
        RECT 114.605 98.845 114.775 99.015 ;
        RECT 115.065 98.845 115.235 99.015 ;
        RECT 115.525 98.845 115.695 99.015 ;
        RECT 115.985 98.845 116.155 99.015 ;
        RECT 116.445 98.845 116.615 99.015 ;
        RECT 116.905 98.845 117.075 99.015 ;
        RECT 117.365 98.845 117.535 99.015 ;
        RECT 117.825 98.845 117.995 99.015 ;
        RECT 118.285 98.845 118.455 99.015 ;
        RECT 118.745 98.845 118.915 99.015 ;
        RECT 119.205 98.845 119.375 99.015 ;
        RECT 119.665 98.845 119.835 99.015 ;
        RECT 120.125 98.845 120.295 99.015 ;
        RECT 120.585 98.845 120.755 99.015 ;
        RECT 121.045 98.845 121.215 99.015 ;
        RECT 121.505 98.845 121.675 99.015 ;
        RECT 121.965 98.845 122.135 99.015 ;
        RECT 122.425 98.845 122.595 99.015 ;
        RECT 122.885 98.845 123.055 99.015 ;
        RECT 123.345 98.845 123.515 99.015 ;
        RECT 123.805 98.845 123.975 99.015 ;
        RECT 124.265 98.845 124.435 99.015 ;
        RECT 124.725 98.845 124.895 99.015 ;
        RECT 125.185 98.845 125.355 99.015 ;
        RECT 125.645 98.845 125.815 99.015 ;
        RECT 126.105 98.845 126.275 99.015 ;
        RECT 126.565 98.845 126.735 99.015 ;
        RECT 127.025 98.845 127.195 99.015 ;
        RECT 127.485 98.845 127.655 99.015 ;
        RECT 127.945 98.845 128.115 99.015 ;
        RECT 128.405 98.845 128.575 99.015 ;
        RECT 128.865 98.845 129.035 99.015 ;
        RECT 129.325 98.845 129.495 99.015 ;
        RECT 129.785 98.845 129.955 99.015 ;
        RECT 130.245 98.845 130.415 99.015 ;
        RECT 130.705 98.845 130.875 99.015 ;
        RECT 131.165 98.845 131.335 99.015 ;
        RECT 131.625 98.845 131.795 99.015 ;
        RECT 132.085 98.845 132.255 99.015 ;
        RECT 132.545 98.845 132.715 99.015 ;
        RECT 133.005 98.845 133.175 99.015 ;
        RECT 133.465 98.845 133.635 99.015 ;
        RECT 133.925 98.845 134.095 99.015 ;
        RECT 134.385 98.845 134.555 99.015 ;
        RECT 134.845 98.845 135.015 99.015 ;
        RECT 135.305 98.845 135.475 99.015 ;
        RECT 135.765 98.845 135.935 99.015 ;
        RECT 136.225 98.845 136.395 99.015 ;
        RECT 136.685 98.845 136.855 99.015 ;
        RECT 137.145 98.845 137.315 99.015 ;
        RECT 137.605 98.845 137.775 99.015 ;
        RECT 138.065 98.845 138.235 99.015 ;
        RECT 138.525 98.845 138.695 99.015 ;
        RECT 138.985 98.845 139.155 99.015 ;
        RECT 61.705 98.335 61.875 98.505 ;
        RECT 60.785 97.655 60.955 97.825 ;
        RECT 50.665 96.125 50.835 96.295 ;
        RECT 51.125 96.125 51.295 96.295 ;
        RECT 51.585 96.125 51.755 96.295 ;
        RECT 52.045 96.125 52.215 96.295 ;
        RECT 52.505 96.125 52.675 96.295 ;
        RECT 52.965 96.125 53.135 96.295 ;
        RECT 53.425 96.125 53.595 96.295 ;
        RECT 53.885 96.125 54.055 96.295 ;
        RECT 54.345 96.125 54.515 96.295 ;
        RECT 54.805 96.125 54.975 96.295 ;
        RECT 55.265 96.125 55.435 96.295 ;
        RECT 55.725 96.125 55.895 96.295 ;
        RECT 56.185 96.125 56.355 96.295 ;
        RECT 56.645 96.125 56.815 96.295 ;
        RECT 57.105 96.125 57.275 96.295 ;
        RECT 57.565 96.125 57.735 96.295 ;
        RECT 58.025 96.125 58.195 96.295 ;
        RECT 58.485 96.125 58.655 96.295 ;
        RECT 58.945 96.125 59.115 96.295 ;
        RECT 59.405 96.125 59.575 96.295 ;
        RECT 59.865 96.125 60.035 96.295 ;
        RECT 60.325 96.125 60.495 96.295 ;
        RECT 60.785 96.125 60.955 96.295 ;
        RECT 61.245 96.125 61.415 96.295 ;
        RECT 61.705 96.125 61.875 96.295 ;
        RECT 62.165 96.125 62.335 96.295 ;
        RECT 62.625 96.125 62.795 96.295 ;
        RECT 63.085 96.125 63.255 96.295 ;
        RECT 63.545 96.125 63.715 96.295 ;
        RECT 64.005 96.125 64.175 96.295 ;
        RECT 64.465 96.125 64.635 96.295 ;
        RECT 64.925 96.125 65.095 96.295 ;
        RECT 65.385 96.125 65.555 96.295 ;
        RECT 65.845 96.125 66.015 96.295 ;
        RECT 66.305 96.125 66.475 96.295 ;
        RECT 66.765 96.125 66.935 96.295 ;
        RECT 67.225 96.125 67.395 96.295 ;
        RECT 67.685 96.125 67.855 96.295 ;
        RECT 68.145 96.125 68.315 96.295 ;
        RECT 68.605 96.125 68.775 96.295 ;
        RECT 69.065 96.125 69.235 96.295 ;
        RECT 69.525 96.125 69.695 96.295 ;
        RECT 69.985 96.125 70.155 96.295 ;
        RECT 70.445 96.125 70.615 96.295 ;
        RECT 70.905 96.125 71.075 96.295 ;
        RECT 71.365 96.125 71.535 96.295 ;
        RECT 71.825 96.125 71.995 96.295 ;
        RECT 72.285 96.125 72.455 96.295 ;
        RECT 72.745 96.125 72.915 96.295 ;
        RECT 73.205 96.125 73.375 96.295 ;
        RECT 73.665 96.125 73.835 96.295 ;
        RECT 74.125 96.125 74.295 96.295 ;
        RECT 74.585 96.125 74.755 96.295 ;
        RECT 75.045 96.125 75.215 96.295 ;
        RECT 75.505 96.125 75.675 96.295 ;
        RECT 75.965 96.125 76.135 96.295 ;
        RECT 76.425 96.125 76.595 96.295 ;
        RECT 76.885 96.125 77.055 96.295 ;
        RECT 77.345 96.125 77.515 96.295 ;
        RECT 77.805 96.125 77.975 96.295 ;
        RECT 78.265 96.125 78.435 96.295 ;
        RECT 78.725 96.125 78.895 96.295 ;
        RECT 79.185 96.125 79.355 96.295 ;
        RECT 79.645 96.125 79.815 96.295 ;
        RECT 80.105 96.125 80.275 96.295 ;
        RECT 80.565 96.125 80.735 96.295 ;
        RECT 81.025 96.125 81.195 96.295 ;
        RECT 81.485 96.125 81.655 96.295 ;
        RECT 81.945 96.125 82.115 96.295 ;
        RECT 82.405 96.125 82.575 96.295 ;
        RECT 82.865 96.125 83.035 96.295 ;
        RECT 83.325 96.125 83.495 96.295 ;
        RECT 83.785 96.125 83.955 96.295 ;
        RECT 84.245 96.125 84.415 96.295 ;
        RECT 84.705 96.125 84.875 96.295 ;
        RECT 85.165 96.125 85.335 96.295 ;
        RECT 85.625 96.125 85.795 96.295 ;
        RECT 86.085 96.125 86.255 96.295 ;
        RECT 86.545 96.125 86.715 96.295 ;
        RECT 87.005 96.125 87.175 96.295 ;
        RECT 87.465 96.125 87.635 96.295 ;
        RECT 87.925 96.125 88.095 96.295 ;
        RECT 88.385 96.125 88.555 96.295 ;
        RECT 88.845 96.125 89.015 96.295 ;
        RECT 89.305 96.125 89.475 96.295 ;
        RECT 89.765 96.125 89.935 96.295 ;
        RECT 90.225 96.125 90.395 96.295 ;
        RECT 90.685 96.125 90.855 96.295 ;
        RECT 91.145 96.125 91.315 96.295 ;
        RECT 91.605 96.125 91.775 96.295 ;
        RECT 92.065 96.125 92.235 96.295 ;
        RECT 92.525 96.125 92.695 96.295 ;
        RECT 92.985 96.125 93.155 96.295 ;
        RECT 93.445 96.125 93.615 96.295 ;
        RECT 93.905 96.125 94.075 96.295 ;
        RECT 94.365 96.125 94.535 96.295 ;
        RECT 94.825 96.125 94.995 96.295 ;
        RECT 95.285 96.125 95.455 96.295 ;
        RECT 95.745 96.125 95.915 96.295 ;
        RECT 96.205 96.125 96.375 96.295 ;
        RECT 96.665 96.125 96.835 96.295 ;
        RECT 97.125 96.125 97.295 96.295 ;
        RECT 97.585 96.125 97.755 96.295 ;
        RECT 98.045 96.125 98.215 96.295 ;
        RECT 98.505 96.125 98.675 96.295 ;
        RECT 98.965 96.125 99.135 96.295 ;
        RECT 99.425 96.125 99.595 96.295 ;
        RECT 99.885 96.125 100.055 96.295 ;
        RECT 100.345 96.125 100.515 96.295 ;
        RECT 100.805 96.125 100.975 96.295 ;
        RECT 101.265 96.125 101.435 96.295 ;
        RECT 101.725 96.125 101.895 96.295 ;
        RECT 102.185 96.125 102.355 96.295 ;
        RECT 102.645 96.125 102.815 96.295 ;
        RECT 103.105 96.125 103.275 96.295 ;
        RECT 103.565 96.125 103.735 96.295 ;
        RECT 104.025 96.125 104.195 96.295 ;
        RECT 104.485 96.125 104.655 96.295 ;
        RECT 104.945 96.125 105.115 96.295 ;
        RECT 105.405 96.125 105.575 96.295 ;
        RECT 105.865 96.125 106.035 96.295 ;
        RECT 106.325 96.125 106.495 96.295 ;
        RECT 106.785 96.125 106.955 96.295 ;
        RECT 107.245 96.125 107.415 96.295 ;
        RECT 107.705 96.125 107.875 96.295 ;
        RECT 108.165 96.125 108.335 96.295 ;
        RECT 108.625 96.125 108.795 96.295 ;
        RECT 109.085 96.125 109.255 96.295 ;
        RECT 109.545 96.125 109.715 96.295 ;
        RECT 110.005 96.125 110.175 96.295 ;
        RECT 110.465 96.125 110.635 96.295 ;
        RECT 110.925 96.125 111.095 96.295 ;
        RECT 111.385 96.125 111.555 96.295 ;
        RECT 111.845 96.125 112.015 96.295 ;
        RECT 112.305 96.125 112.475 96.295 ;
        RECT 112.765 96.125 112.935 96.295 ;
        RECT 113.225 96.125 113.395 96.295 ;
        RECT 113.685 96.125 113.855 96.295 ;
        RECT 114.145 96.125 114.315 96.295 ;
        RECT 114.605 96.125 114.775 96.295 ;
        RECT 115.065 96.125 115.235 96.295 ;
        RECT 115.525 96.125 115.695 96.295 ;
        RECT 115.985 96.125 116.155 96.295 ;
        RECT 116.445 96.125 116.615 96.295 ;
        RECT 116.905 96.125 117.075 96.295 ;
        RECT 117.365 96.125 117.535 96.295 ;
        RECT 117.825 96.125 117.995 96.295 ;
        RECT 118.285 96.125 118.455 96.295 ;
        RECT 118.745 96.125 118.915 96.295 ;
        RECT 119.205 96.125 119.375 96.295 ;
        RECT 119.665 96.125 119.835 96.295 ;
        RECT 120.125 96.125 120.295 96.295 ;
        RECT 120.585 96.125 120.755 96.295 ;
        RECT 121.045 96.125 121.215 96.295 ;
        RECT 121.505 96.125 121.675 96.295 ;
        RECT 121.965 96.125 122.135 96.295 ;
        RECT 122.425 96.125 122.595 96.295 ;
        RECT 122.885 96.125 123.055 96.295 ;
        RECT 123.345 96.125 123.515 96.295 ;
        RECT 123.805 96.125 123.975 96.295 ;
        RECT 124.265 96.125 124.435 96.295 ;
        RECT 124.725 96.125 124.895 96.295 ;
        RECT 125.185 96.125 125.355 96.295 ;
        RECT 125.645 96.125 125.815 96.295 ;
        RECT 126.105 96.125 126.275 96.295 ;
        RECT 126.565 96.125 126.735 96.295 ;
        RECT 127.025 96.125 127.195 96.295 ;
        RECT 127.485 96.125 127.655 96.295 ;
        RECT 127.945 96.125 128.115 96.295 ;
        RECT 128.405 96.125 128.575 96.295 ;
        RECT 128.865 96.125 129.035 96.295 ;
        RECT 129.325 96.125 129.495 96.295 ;
        RECT 129.785 96.125 129.955 96.295 ;
        RECT 130.245 96.125 130.415 96.295 ;
        RECT 130.705 96.125 130.875 96.295 ;
        RECT 131.165 96.125 131.335 96.295 ;
        RECT 131.625 96.125 131.795 96.295 ;
        RECT 132.085 96.125 132.255 96.295 ;
        RECT 132.545 96.125 132.715 96.295 ;
        RECT 133.005 96.125 133.175 96.295 ;
        RECT 133.465 96.125 133.635 96.295 ;
        RECT 133.925 96.125 134.095 96.295 ;
        RECT 134.385 96.125 134.555 96.295 ;
        RECT 134.845 96.125 135.015 96.295 ;
        RECT 135.305 96.125 135.475 96.295 ;
        RECT 135.765 96.125 135.935 96.295 ;
        RECT 136.225 96.125 136.395 96.295 ;
        RECT 136.685 96.125 136.855 96.295 ;
        RECT 137.145 96.125 137.315 96.295 ;
        RECT 137.605 96.125 137.775 96.295 ;
        RECT 138.065 96.125 138.235 96.295 ;
        RECT 138.525 96.125 138.695 96.295 ;
        RECT 138.985 96.125 139.155 96.295 ;
        RECT 61.705 94.595 61.875 94.765 ;
        RECT 62.625 94.595 62.795 94.765 ;
        RECT 61.705 93.915 61.875 94.085 ;
        RECT 50.665 93.405 50.835 93.575 ;
        RECT 51.125 93.405 51.295 93.575 ;
        RECT 51.585 93.405 51.755 93.575 ;
        RECT 52.045 93.405 52.215 93.575 ;
        RECT 52.505 93.405 52.675 93.575 ;
        RECT 52.965 93.405 53.135 93.575 ;
        RECT 53.425 93.405 53.595 93.575 ;
        RECT 53.885 93.405 54.055 93.575 ;
        RECT 54.345 93.405 54.515 93.575 ;
        RECT 54.805 93.405 54.975 93.575 ;
        RECT 55.265 93.405 55.435 93.575 ;
        RECT 55.725 93.405 55.895 93.575 ;
        RECT 56.185 93.405 56.355 93.575 ;
        RECT 56.645 93.405 56.815 93.575 ;
        RECT 57.105 93.405 57.275 93.575 ;
        RECT 57.565 93.405 57.735 93.575 ;
        RECT 58.025 93.405 58.195 93.575 ;
        RECT 58.485 93.405 58.655 93.575 ;
        RECT 58.945 93.405 59.115 93.575 ;
        RECT 59.405 93.405 59.575 93.575 ;
        RECT 59.865 93.405 60.035 93.575 ;
        RECT 60.325 93.405 60.495 93.575 ;
        RECT 60.785 93.405 60.955 93.575 ;
        RECT 61.245 93.405 61.415 93.575 ;
        RECT 61.705 93.405 61.875 93.575 ;
        RECT 62.165 93.405 62.335 93.575 ;
        RECT 62.625 93.405 62.795 93.575 ;
        RECT 63.085 93.405 63.255 93.575 ;
        RECT 63.545 93.405 63.715 93.575 ;
        RECT 64.005 93.405 64.175 93.575 ;
        RECT 64.465 93.405 64.635 93.575 ;
        RECT 64.925 93.405 65.095 93.575 ;
        RECT 65.385 93.405 65.555 93.575 ;
        RECT 65.845 93.405 66.015 93.575 ;
        RECT 66.305 93.405 66.475 93.575 ;
        RECT 66.765 93.405 66.935 93.575 ;
        RECT 67.225 93.405 67.395 93.575 ;
        RECT 67.685 93.405 67.855 93.575 ;
        RECT 68.145 93.405 68.315 93.575 ;
        RECT 68.605 93.405 68.775 93.575 ;
        RECT 69.065 93.405 69.235 93.575 ;
        RECT 69.525 93.405 69.695 93.575 ;
        RECT 69.985 93.405 70.155 93.575 ;
        RECT 70.445 93.405 70.615 93.575 ;
        RECT 70.905 93.405 71.075 93.575 ;
        RECT 71.365 93.405 71.535 93.575 ;
        RECT 71.825 93.405 71.995 93.575 ;
        RECT 72.285 93.405 72.455 93.575 ;
        RECT 72.745 93.405 72.915 93.575 ;
        RECT 73.205 93.405 73.375 93.575 ;
        RECT 73.665 93.405 73.835 93.575 ;
        RECT 74.125 93.405 74.295 93.575 ;
        RECT 74.585 93.405 74.755 93.575 ;
        RECT 75.045 93.405 75.215 93.575 ;
        RECT 75.505 93.405 75.675 93.575 ;
        RECT 75.965 93.405 76.135 93.575 ;
        RECT 76.425 93.405 76.595 93.575 ;
        RECT 76.885 93.405 77.055 93.575 ;
        RECT 77.345 93.405 77.515 93.575 ;
        RECT 77.805 93.405 77.975 93.575 ;
        RECT 78.265 93.405 78.435 93.575 ;
        RECT 78.725 93.405 78.895 93.575 ;
        RECT 79.185 93.405 79.355 93.575 ;
        RECT 79.645 93.405 79.815 93.575 ;
        RECT 80.105 93.405 80.275 93.575 ;
        RECT 80.565 93.405 80.735 93.575 ;
        RECT 81.025 93.405 81.195 93.575 ;
        RECT 81.485 93.405 81.655 93.575 ;
        RECT 81.945 93.405 82.115 93.575 ;
        RECT 82.405 93.405 82.575 93.575 ;
        RECT 82.865 93.405 83.035 93.575 ;
        RECT 83.325 93.405 83.495 93.575 ;
        RECT 83.785 93.405 83.955 93.575 ;
        RECT 84.245 93.405 84.415 93.575 ;
        RECT 84.705 93.405 84.875 93.575 ;
        RECT 85.165 93.405 85.335 93.575 ;
        RECT 85.625 93.405 85.795 93.575 ;
        RECT 86.085 93.405 86.255 93.575 ;
        RECT 86.545 93.405 86.715 93.575 ;
        RECT 87.005 93.405 87.175 93.575 ;
        RECT 87.465 93.405 87.635 93.575 ;
        RECT 87.925 93.405 88.095 93.575 ;
        RECT 88.385 93.405 88.555 93.575 ;
        RECT 88.845 93.405 89.015 93.575 ;
        RECT 89.305 93.405 89.475 93.575 ;
        RECT 89.765 93.405 89.935 93.575 ;
        RECT 90.225 93.405 90.395 93.575 ;
        RECT 90.685 93.405 90.855 93.575 ;
        RECT 91.145 93.405 91.315 93.575 ;
        RECT 91.605 93.405 91.775 93.575 ;
        RECT 92.065 93.405 92.235 93.575 ;
        RECT 92.525 93.405 92.695 93.575 ;
        RECT 92.985 93.405 93.155 93.575 ;
        RECT 93.445 93.405 93.615 93.575 ;
        RECT 93.905 93.405 94.075 93.575 ;
        RECT 94.365 93.405 94.535 93.575 ;
        RECT 94.825 93.405 94.995 93.575 ;
        RECT 95.285 93.405 95.455 93.575 ;
        RECT 95.745 93.405 95.915 93.575 ;
        RECT 96.205 93.405 96.375 93.575 ;
        RECT 96.665 93.405 96.835 93.575 ;
        RECT 97.125 93.405 97.295 93.575 ;
        RECT 97.585 93.405 97.755 93.575 ;
        RECT 98.045 93.405 98.215 93.575 ;
        RECT 98.505 93.405 98.675 93.575 ;
        RECT 98.965 93.405 99.135 93.575 ;
        RECT 99.425 93.405 99.595 93.575 ;
        RECT 99.885 93.405 100.055 93.575 ;
        RECT 100.345 93.405 100.515 93.575 ;
        RECT 100.805 93.405 100.975 93.575 ;
        RECT 101.265 93.405 101.435 93.575 ;
        RECT 101.725 93.405 101.895 93.575 ;
        RECT 102.185 93.405 102.355 93.575 ;
        RECT 102.645 93.405 102.815 93.575 ;
        RECT 103.105 93.405 103.275 93.575 ;
        RECT 103.565 93.405 103.735 93.575 ;
        RECT 104.025 93.405 104.195 93.575 ;
        RECT 104.485 93.405 104.655 93.575 ;
        RECT 104.945 93.405 105.115 93.575 ;
        RECT 105.405 93.405 105.575 93.575 ;
        RECT 105.865 93.405 106.035 93.575 ;
        RECT 106.325 93.405 106.495 93.575 ;
        RECT 106.785 93.405 106.955 93.575 ;
        RECT 107.245 93.405 107.415 93.575 ;
        RECT 107.705 93.405 107.875 93.575 ;
        RECT 108.165 93.405 108.335 93.575 ;
        RECT 108.625 93.405 108.795 93.575 ;
        RECT 109.085 93.405 109.255 93.575 ;
        RECT 109.545 93.405 109.715 93.575 ;
        RECT 110.005 93.405 110.175 93.575 ;
        RECT 110.465 93.405 110.635 93.575 ;
        RECT 110.925 93.405 111.095 93.575 ;
        RECT 111.385 93.405 111.555 93.575 ;
        RECT 111.845 93.405 112.015 93.575 ;
        RECT 112.305 93.405 112.475 93.575 ;
        RECT 112.765 93.405 112.935 93.575 ;
        RECT 113.225 93.405 113.395 93.575 ;
        RECT 113.685 93.405 113.855 93.575 ;
        RECT 114.145 93.405 114.315 93.575 ;
        RECT 114.605 93.405 114.775 93.575 ;
        RECT 115.065 93.405 115.235 93.575 ;
        RECT 115.525 93.405 115.695 93.575 ;
        RECT 115.985 93.405 116.155 93.575 ;
        RECT 116.445 93.405 116.615 93.575 ;
        RECT 116.905 93.405 117.075 93.575 ;
        RECT 117.365 93.405 117.535 93.575 ;
        RECT 117.825 93.405 117.995 93.575 ;
        RECT 118.285 93.405 118.455 93.575 ;
        RECT 118.745 93.405 118.915 93.575 ;
        RECT 119.205 93.405 119.375 93.575 ;
        RECT 119.665 93.405 119.835 93.575 ;
        RECT 120.125 93.405 120.295 93.575 ;
        RECT 120.585 93.405 120.755 93.575 ;
        RECT 121.045 93.405 121.215 93.575 ;
        RECT 121.505 93.405 121.675 93.575 ;
        RECT 121.965 93.405 122.135 93.575 ;
        RECT 122.425 93.405 122.595 93.575 ;
        RECT 122.885 93.405 123.055 93.575 ;
        RECT 123.345 93.405 123.515 93.575 ;
        RECT 123.805 93.405 123.975 93.575 ;
        RECT 124.265 93.405 124.435 93.575 ;
        RECT 124.725 93.405 124.895 93.575 ;
        RECT 125.185 93.405 125.355 93.575 ;
        RECT 125.645 93.405 125.815 93.575 ;
        RECT 126.105 93.405 126.275 93.575 ;
        RECT 126.565 93.405 126.735 93.575 ;
        RECT 127.025 93.405 127.195 93.575 ;
        RECT 127.485 93.405 127.655 93.575 ;
        RECT 127.945 93.405 128.115 93.575 ;
        RECT 128.405 93.405 128.575 93.575 ;
        RECT 128.865 93.405 129.035 93.575 ;
        RECT 129.325 93.405 129.495 93.575 ;
        RECT 129.785 93.405 129.955 93.575 ;
        RECT 130.245 93.405 130.415 93.575 ;
        RECT 130.705 93.405 130.875 93.575 ;
        RECT 131.165 93.405 131.335 93.575 ;
        RECT 131.625 93.405 131.795 93.575 ;
        RECT 132.085 93.405 132.255 93.575 ;
        RECT 132.545 93.405 132.715 93.575 ;
        RECT 133.005 93.405 133.175 93.575 ;
        RECT 133.465 93.405 133.635 93.575 ;
        RECT 133.925 93.405 134.095 93.575 ;
        RECT 134.385 93.405 134.555 93.575 ;
        RECT 134.845 93.405 135.015 93.575 ;
        RECT 135.305 93.405 135.475 93.575 ;
        RECT 135.765 93.405 135.935 93.575 ;
        RECT 136.225 93.405 136.395 93.575 ;
        RECT 136.685 93.405 136.855 93.575 ;
        RECT 137.145 93.405 137.315 93.575 ;
        RECT 137.605 93.405 137.775 93.575 ;
        RECT 138.065 93.405 138.235 93.575 ;
        RECT 138.525 93.405 138.695 93.575 ;
        RECT 138.985 93.405 139.155 93.575 ;
        RECT 58.025 92.895 58.195 93.065 ;
        RECT 57.565 91.875 57.735 92.045 ;
        RECT 58.485 92.895 58.655 93.065 ;
        RECT 60.325 91.195 60.495 91.365 ;
        RECT 60.785 92.895 60.955 93.065 ;
        RECT 63.085 92.555 63.255 92.725 ;
        RECT 63.545 91.875 63.715 92.045 ;
        RECT 64.925 92.215 65.095 92.385 ;
        RECT 66.765 92.555 66.935 92.725 ;
        RECT 66.305 92.215 66.475 92.385 ;
        RECT 50.665 90.685 50.835 90.855 ;
        RECT 51.125 90.685 51.295 90.855 ;
        RECT 51.585 90.685 51.755 90.855 ;
        RECT 52.045 90.685 52.215 90.855 ;
        RECT 52.505 90.685 52.675 90.855 ;
        RECT 52.965 90.685 53.135 90.855 ;
        RECT 53.425 90.685 53.595 90.855 ;
        RECT 53.885 90.685 54.055 90.855 ;
        RECT 54.345 90.685 54.515 90.855 ;
        RECT 54.805 90.685 54.975 90.855 ;
        RECT 55.265 90.685 55.435 90.855 ;
        RECT 55.725 90.685 55.895 90.855 ;
        RECT 56.185 90.685 56.355 90.855 ;
        RECT 56.645 90.685 56.815 90.855 ;
        RECT 57.105 90.685 57.275 90.855 ;
        RECT 57.565 90.685 57.735 90.855 ;
        RECT 58.025 90.685 58.195 90.855 ;
        RECT 58.485 90.685 58.655 90.855 ;
        RECT 58.945 90.685 59.115 90.855 ;
        RECT 59.405 90.685 59.575 90.855 ;
        RECT 59.865 90.685 60.035 90.855 ;
        RECT 60.325 90.685 60.495 90.855 ;
        RECT 60.785 90.685 60.955 90.855 ;
        RECT 61.245 90.685 61.415 90.855 ;
        RECT 61.705 90.685 61.875 90.855 ;
        RECT 62.165 90.685 62.335 90.855 ;
        RECT 62.625 90.685 62.795 90.855 ;
        RECT 63.085 90.685 63.255 90.855 ;
        RECT 63.545 90.685 63.715 90.855 ;
        RECT 64.005 90.685 64.175 90.855 ;
        RECT 64.465 90.685 64.635 90.855 ;
        RECT 64.925 90.685 65.095 90.855 ;
        RECT 65.385 90.685 65.555 90.855 ;
        RECT 65.845 90.685 66.015 90.855 ;
        RECT 66.305 90.685 66.475 90.855 ;
        RECT 66.765 90.685 66.935 90.855 ;
        RECT 67.225 90.685 67.395 90.855 ;
        RECT 67.685 90.685 67.855 90.855 ;
        RECT 68.145 90.685 68.315 90.855 ;
        RECT 68.605 90.685 68.775 90.855 ;
        RECT 69.065 90.685 69.235 90.855 ;
        RECT 69.525 90.685 69.695 90.855 ;
        RECT 69.985 90.685 70.155 90.855 ;
        RECT 70.445 90.685 70.615 90.855 ;
        RECT 70.905 90.685 71.075 90.855 ;
        RECT 71.365 90.685 71.535 90.855 ;
        RECT 71.825 90.685 71.995 90.855 ;
        RECT 72.285 90.685 72.455 90.855 ;
        RECT 72.745 90.685 72.915 90.855 ;
        RECT 73.205 90.685 73.375 90.855 ;
        RECT 73.665 90.685 73.835 90.855 ;
        RECT 74.125 90.685 74.295 90.855 ;
        RECT 74.585 90.685 74.755 90.855 ;
        RECT 75.045 90.685 75.215 90.855 ;
        RECT 75.505 90.685 75.675 90.855 ;
        RECT 75.965 90.685 76.135 90.855 ;
        RECT 76.425 90.685 76.595 90.855 ;
        RECT 76.885 90.685 77.055 90.855 ;
        RECT 77.345 90.685 77.515 90.855 ;
        RECT 77.805 90.685 77.975 90.855 ;
        RECT 78.265 90.685 78.435 90.855 ;
        RECT 78.725 90.685 78.895 90.855 ;
        RECT 79.185 90.685 79.355 90.855 ;
        RECT 79.645 90.685 79.815 90.855 ;
        RECT 80.105 90.685 80.275 90.855 ;
        RECT 80.565 90.685 80.735 90.855 ;
        RECT 81.025 90.685 81.195 90.855 ;
        RECT 81.485 90.685 81.655 90.855 ;
        RECT 81.945 90.685 82.115 90.855 ;
        RECT 82.405 90.685 82.575 90.855 ;
        RECT 82.865 90.685 83.035 90.855 ;
        RECT 83.325 90.685 83.495 90.855 ;
        RECT 83.785 90.685 83.955 90.855 ;
        RECT 84.245 90.685 84.415 90.855 ;
        RECT 84.705 90.685 84.875 90.855 ;
        RECT 85.165 90.685 85.335 90.855 ;
        RECT 85.625 90.685 85.795 90.855 ;
        RECT 86.085 90.685 86.255 90.855 ;
        RECT 86.545 90.685 86.715 90.855 ;
        RECT 87.005 90.685 87.175 90.855 ;
        RECT 87.465 90.685 87.635 90.855 ;
        RECT 87.925 90.685 88.095 90.855 ;
        RECT 88.385 90.685 88.555 90.855 ;
        RECT 88.845 90.685 89.015 90.855 ;
        RECT 89.305 90.685 89.475 90.855 ;
        RECT 89.765 90.685 89.935 90.855 ;
        RECT 90.225 90.685 90.395 90.855 ;
        RECT 90.685 90.685 90.855 90.855 ;
        RECT 91.145 90.685 91.315 90.855 ;
        RECT 91.605 90.685 91.775 90.855 ;
        RECT 92.065 90.685 92.235 90.855 ;
        RECT 92.525 90.685 92.695 90.855 ;
        RECT 92.985 90.685 93.155 90.855 ;
        RECT 93.445 90.685 93.615 90.855 ;
        RECT 93.905 90.685 94.075 90.855 ;
        RECT 94.365 90.685 94.535 90.855 ;
        RECT 94.825 90.685 94.995 90.855 ;
        RECT 95.285 90.685 95.455 90.855 ;
        RECT 95.745 90.685 95.915 90.855 ;
        RECT 96.205 90.685 96.375 90.855 ;
        RECT 96.665 90.685 96.835 90.855 ;
        RECT 97.125 90.685 97.295 90.855 ;
        RECT 97.585 90.685 97.755 90.855 ;
        RECT 98.045 90.685 98.215 90.855 ;
        RECT 98.505 90.685 98.675 90.855 ;
        RECT 98.965 90.685 99.135 90.855 ;
        RECT 99.425 90.685 99.595 90.855 ;
        RECT 99.885 90.685 100.055 90.855 ;
        RECT 100.345 90.685 100.515 90.855 ;
        RECT 100.805 90.685 100.975 90.855 ;
        RECT 101.265 90.685 101.435 90.855 ;
        RECT 101.725 90.685 101.895 90.855 ;
        RECT 102.185 90.685 102.355 90.855 ;
        RECT 102.645 90.685 102.815 90.855 ;
        RECT 103.105 90.685 103.275 90.855 ;
        RECT 103.565 90.685 103.735 90.855 ;
        RECT 104.025 90.685 104.195 90.855 ;
        RECT 104.485 90.685 104.655 90.855 ;
        RECT 104.945 90.685 105.115 90.855 ;
        RECT 105.405 90.685 105.575 90.855 ;
        RECT 105.865 90.685 106.035 90.855 ;
        RECT 106.325 90.685 106.495 90.855 ;
        RECT 106.785 90.685 106.955 90.855 ;
        RECT 107.245 90.685 107.415 90.855 ;
        RECT 107.705 90.685 107.875 90.855 ;
        RECT 108.165 90.685 108.335 90.855 ;
        RECT 108.625 90.685 108.795 90.855 ;
        RECT 109.085 90.685 109.255 90.855 ;
        RECT 109.545 90.685 109.715 90.855 ;
        RECT 110.005 90.685 110.175 90.855 ;
        RECT 110.465 90.685 110.635 90.855 ;
        RECT 110.925 90.685 111.095 90.855 ;
        RECT 111.385 90.685 111.555 90.855 ;
        RECT 111.845 90.685 112.015 90.855 ;
        RECT 112.305 90.685 112.475 90.855 ;
        RECT 112.765 90.685 112.935 90.855 ;
        RECT 113.225 90.685 113.395 90.855 ;
        RECT 113.685 90.685 113.855 90.855 ;
        RECT 114.145 90.685 114.315 90.855 ;
        RECT 114.605 90.685 114.775 90.855 ;
        RECT 115.065 90.685 115.235 90.855 ;
        RECT 115.525 90.685 115.695 90.855 ;
        RECT 115.985 90.685 116.155 90.855 ;
        RECT 116.445 90.685 116.615 90.855 ;
        RECT 116.905 90.685 117.075 90.855 ;
        RECT 117.365 90.685 117.535 90.855 ;
        RECT 117.825 90.685 117.995 90.855 ;
        RECT 118.285 90.685 118.455 90.855 ;
        RECT 118.745 90.685 118.915 90.855 ;
        RECT 119.205 90.685 119.375 90.855 ;
        RECT 119.665 90.685 119.835 90.855 ;
        RECT 120.125 90.685 120.295 90.855 ;
        RECT 120.585 90.685 120.755 90.855 ;
        RECT 121.045 90.685 121.215 90.855 ;
        RECT 121.505 90.685 121.675 90.855 ;
        RECT 121.965 90.685 122.135 90.855 ;
        RECT 122.425 90.685 122.595 90.855 ;
        RECT 122.885 90.685 123.055 90.855 ;
        RECT 123.345 90.685 123.515 90.855 ;
        RECT 123.805 90.685 123.975 90.855 ;
        RECT 124.265 90.685 124.435 90.855 ;
        RECT 124.725 90.685 124.895 90.855 ;
        RECT 125.185 90.685 125.355 90.855 ;
        RECT 125.645 90.685 125.815 90.855 ;
        RECT 126.105 90.685 126.275 90.855 ;
        RECT 126.565 90.685 126.735 90.855 ;
        RECT 127.025 90.685 127.195 90.855 ;
        RECT 127.485 90.685 127.655 90.855 ;
        RECT 127.945 90.685 128.115 90.855 ;
        RECT 128.405 90.685 128.575 90.855 ;
        RECT 128.865 90.685 129.035 90.855 ;
        RECT 129.325 90.685 129.495 90.855 ;
        RECT 129.785 90.685 129.955 90.855 ;
        RECT 130.245 90.685 130.415 90.855 ;
        RECT 130.705 90.685 130.875 90.855 ;
        RECT 131.165 90.685 131.335 90.855 ;
        RECT 131.625 90.685 131.795 90.855 ;
        RECT 132.085 90.685 132.255 90.855 ;
        RECT 132.545 90.685 132.715 90.855 ;
        RECT 133.005 90.685 133.175 90.855 ;
        RECT 133.465 90.685 133.635 90.855 ;
        RECT 133.925 90.685 134.095 90.855 ;
        RECT 134.385 90.685 134.555 90.855 ;
        RECT 134.845 90.685 135.015 90.855 ;
        RECT 135.305 90.685 135.475 90.855 ;
        RECT 135.765 90.685 135.935 90.855 ;
        RECT 136.225 90.685 136.395 90.855 ;
        RECT 136.685 90.685 136.855 90.855 ;
        RECT 137.145 90.685 137.315 90.855 ;
        RECT 137.605 90.685 137.775 90.855 ;
        RECT 138.065 90.685 138.235 90.855 ;
        RECT 138.525 90.685 138.695 90.855 ;
        RECT 138.985 90.685 139.155 90.855 ;
        RECT 60.325 89.155 60.495 89.325 ;
        RECT 62.165 90.175 62.335 90.345 ;
        RECT 61.705 89.155 61.875 89.325 ;
        RECT 50.665 87.965 50.835 88.135 ;
        RECT 51.125 87.965 51.295 88.135 ;
        RECT 51.585 87.965 51.755 88.135 ;
        RECT 52.045 87.965 52.215 88.135 ;
        RECT 52.505 87.965 52.675 88.135 ;
        RECT 52.965 87.965 53.135 88.135 ;
        RECT 53.425 87.965 53.595 88.135 ;
        RECT 53.885 87.965 54.055 88.135 ;
        RECT 54.345 87.965 54.515 88.135 ;
        RECT 54.805 87.965 54.975 88.135 ;
        RECT 55.265 87.965 55.435 88.135 ;
        RECT 55.725 87.965 55.895 88.135 ;
        RECT 56.185 87.965 56.355 88.135 ;
        RECT 56.645 87.965 56.815 88.135 ;
        RECT 57.105 87.965 57.275 88.135 ;
        RECT 57.565 87.965 57.735 88.135 ;
        RECT 58.025 87.965 58.195 88.135 ;
        RECT 58.485 87.965 58.655 88.135 ;
        RECT 58.945 87.965 59.115 88.135 ;
        RECT 59.405 87.965 59.575 88.135 ;
        RECT 59.865 87.965 60.035 88.135 ;
        RECT 60.325 87.965 60.495 88.135 ;
        RECT 60.785 87.965 60.955 88.135 ;
        RECT 61.245 87.965 61.415 88.135 ;
        RECT 61.705 87.965 61.875 88.135 ;
        RECT 62.165 87.965 62.335 88.135 ;
        RECT 62.625 87.965 62.795 88.135 ;
        RECT 63.085 87.965 63.255 88.135 ;
        RECT 63.545 87.965 63.715 88.135 ;
        RECT 64.005 87.965 64.175 88.135 ;
        RECT 64.465 87.965 64.635 88.135 ;
        RECT 64.925 87.965 65.095 88.135 ;
        RECT 65.385 87.965 65.555 88.135 ;
        RECT 65.845 87.965 66.015 88.135 ;
        RECT 66.305 87.965 66.475 88.135 ;
        RECT 66.765 87.965 66.935 88.135 ;
        RECT 67.225 87.965 67.395 88.135 ;
        RECT 67.685 87.965 67.855 88.135 ;
        RECT 68.145 87.965 68.315 88.135 ;
        RECT 68.605 87.965 68.775 88.135 ;
        RECT 69.065 87.965 69.235 88.135 ;
        RECT 69.525 87.965 69.695 88.135 ;
        RECT 69.985 87.965 70.155 88.135 ;
        RECT 70.445 87.965 70.615 88.135 ;
        RECT 70.905 87.965 71.075 88.135 ;
        RECT 71.365 87.965 71.535 88.135 ;
        RECT 71.825 87.965 71.995 88.135 ;
        RECT 72.285 87.965 72.455 88.135 ;
        RECT 72.745 87.965 72.915 88.135 ;
        RECT 73.205 87.965 73.375 88.135 ;
        RECT 73.665 87.965 73.835 88.135 ;
        RECT 74.125 87.965 74.295 88.135 ;
        RECT 74.585 87.965 74.755 88.135 ;
        RECT 75.045 87.965 75.215 88.135 ;
        RECT 75.505 87.965 75.675 88.135 ;
        RECT 75.965 87.965 76.135 88.135 ;
        RECT 76.425 87.965 76.595 88.135 ;
        RECT 76.885 87.965 77.055 88.135 ;
        RECT 77.345 87.965 77.515 88.135 ;
        RECT 77.805 87.965 77.975 88.135 ;
        RECT 78.265 87.965 78.435 88.135 ;
        RECT 78.725 87.965 78.895 88.135 ;
        RECT 79.185 87.965 79.355 88.135 ;
        RECT 79.645 87.965 79.815 88.135 ;
        RECT 80.105 87.965 80.275 88.135 ;
        RECT 80.565 87.965 80.735 88.135 ;
        RECT 81.025 87.965 81.195 88.135 ;
        RECT 81.485 87.965 81.655 88.135 ;
        RECT 81.945 87.965 82.115 88.135 ;
        RECT 82.405 87.965 82.575 88.135 ;
        RECT 82.865 87.965 83.035 88.135 ;
        RECT 83.325 87.965 83.495 88.135 ;
        RECT 83.785 87.965 83.955 88.135 ;
        RECT 84.245 87.965 84.415 88.135 ;
        RECT 84.705 87.965 84.875 88.135 ;
        RECT 85.165 87.965 85.335 88.135 ;
        RECT 85.625 87.965 85.795 88.135 ;
        RECT 86.085 87.965 86.255 88.135 ;
        RECT 86.545 87.965 86.715 88.135 ;
        RECT 87.005 87.965 87.175 88.135 ;
        RECT 87.465 87.965 87.635 88.135 ;
        RECT 87.925 87.965 88.095 88.135 ;
        RECT 88.385 87.965 88.555 88.135 ;
        RECT 88.845 87.965 89.015 88.135 ;
        RECT 89.305 87.965 89.475 88.135 ;
        RECT 89.765 87.965 89.935 88.135 ;
        RECT 90.225 87.965 90.395 88.135 ;
        RECT 90.685 87.965 90.855 88.135 ;
        RECT 91.145 87.965 91.315 88.135 ;
        RECT 91.605 87.965 91.775 88.135 ;
        RECT 92.065 87.965 92.235 88.135 ;
        RECT 92.525 87.965 92.695 88.135 ;
        RECT 92.985 87.965 93.155 88.135 ;
        RECT 93.445 87.965 93.615 88.135 ;
        RECT 93.905 87.965 94.075 88.135 ;
        RECT 94.365 87.965 94.535 88.135 ;
        RECT 94.825 87.965 94.995 88.135 ;
        RECT 95.285 87.965 95.455 88.135 ;
        RECT 95.745 87.965 95.915 88.135 ;
        RECT 96.205 87.965 96.375 88.135 ;
        RECT 96.665 87.965 96.835 88.135 ;
        RECT 97.125 87.965 97.295 88.135 ;
        RECT 97.585 87.965 97.755 88.135 ;
        RECT 98.045 87.965 98.215 88.135 ;
        RECT 98.505 87.965 98.675 88.135 ;
        RECT 98.965 87.965 99.135 88.135 ;
        RECT 99.425 87.965 99.595 88.135 ;
        RECT 99.885 87.965 100.055 88.135 ;
        RECT 100.345 87.965 100.515 88.135 ;
        RECT 100.805 87.965 100.975 88.135 ;
        RECT 101.265 87.965 101.435 88.135 ;
        RECT 101.725 87.965 101.895 88.135 ;
        RECT 102.185 87.965 102.355 88.135 ;
        RECT 102.645 87.965 102.815 88.135 ;
        RECT 103.105 87.965 103.275 88.135 ;
        RECT 103.565 87.965 103.735 88.135 ;
        RECT 104.025 87.965 104.195 88.135 ;
        RECT 104.485 87.965 104.655 88.135 ;
        RECT 104.945 87.965 105.115 88.135 ;
        RECT 105.405 87.965 105.575 88.135 ;
        RECT 105.865 87.965 106.035 88.135 ;
        RECT 106.325 87.965 106.495 88.135 ;
        RECT 106.785 87.965 106.955 88.135 ;
        RECT 107.245 87.965 107.415 88.135 ;
        RECT 107.705 87.965 107.875 88.135 ;
        RECT 108.165 87.965 108.335 88.135 ;
        RECT 108.625 87.965 108.795 88.135 ;
        RECT 109.085 87.965 109.255 88.135 ;
        RECT 109.545 87.965 109.715 88.135 ;
        RECT 110.005 87.965 110.175 88.135 ;
        RECT 110.465 87.965 110.635 88.135 ;
        RECT 110.925 87.965 111.095 88.135 ;
        RECT 111.385 87.965 111.555 88.135 ;
        RECT 111.845 87.965 112.015 88.135 ;
        RECT 112.305 87.965 112.475 88.135 ;
        RECT 112.765 87.965 112.935 88.135 ;
        RECT 113.225 87.965 113.395 88.135 ;
        RECT 113.685 87.965 113.855 88.135 ;
        RECT 114.145 87.965 114.315 88.135 ;
        RECT 114.605 87.965 114.775 88.135 ;
        RECT 115.065 87.965 115.235 88.135 ;
        RECT 115.525 87.965 115.695 88.135 ;
        RECT 115.985 87.965 116.155 88.135 ;
        RECT 116.445 87.965 116.615 88.135 ;
        RECT 116.905 87.965 117.075 88.135 ;
        RECT 117.365 87.965 117.535 88.135 ;
        RECT 117.825 87.965 117.995 88.135 ;
        RECT 118.285 87.965 118.455 88.135 ;
        RECT 118.745 87.965 118.915 88.135 ;
        RECT 119.205 87.965 119.375 88.135 ;
        RECT 119.665 87.965 119.835 88.135 ;
        RECT 120.125 87.965 120.295 88.135 ;
        RECT 120.585 87.965 120.755 88.135 ;
        RECT 121.045 87.965 121.215 88.135 ;
        RECT 121.505 87.965 121.675 88.135 ;
        RECT 121.965 87.965 122.135 88.135 ;
        RECT 122.425 87.965 122.595 88.135 ;
        RECT 122.885 87.965 123.055 88.135 ;
        RECT 123.345 87.965 123.515 88.135 ;
        RECT 123.805 87.965 123.975 88.135 ;
        RECT 124.265 87.965 124.435 88.135 ;
        RECT 124.725 87.965 124.895 88.135 ;
        RECT 125.185 87.965 125.355 88.135 ;
        RECT 125.645 87.965 125.815 88.135 ;
        RECT 126.105 87.965 126.275 88.135 ;
        RECT 126.565 87.965 126.735 88.135 ;
        RECT 127.025 87.965 127.195 88.135 ;
        RECT 127.485 87.965 127.655 88.135 ;
        RECT 127.945 87.965 128.115 88.135 ;
        RECT 128.405 87.965 128.575 88.135 ;
        RECT 128.865 87.965 129.035 88.135 ;
        RECT 129.325 87.965 129.495 88.135 ;
        RECT 129.785 87.965 129.955 88.135 ;
        RECT 130.245 87.965 130.415 88.135 ;
        RECT 130.705 87.965 130.875 88.135 ;
        RECT 131.165 87.965 131.335 88.135 ;
        RECT 131.625 87.965 131.795 88.135 ;
        RECT 132.085 87.965 132.255 88.135 ;
        RECT 132.545 87.965 132.715 88.135 ;
        RECT 133.005 87.965 133.175 88.135 ;
        RECT 133.465 87.965 133.635 88.135 ;
        RECT 133.925 87.965 134.095 88.135 ;
        RECT 134.385 87.965 134.555 88.135 ;
        RECT 134.845 87.965 135.015 88.135 ;
        RECT 135.305 87.965 135.475 88.135 ;
        RECT 135.765 87.965 135.935 88.135 ;
        RECT 136.225 87.965 136.395 88.135 ;
        RECT 136.685 87.965 136.855 88.135 ;
        RECT 137.145 87.965 137.315 88.135 ;
        RECT 137.605 87.965 137.775 88.135 ;
        RECT 138.065 87.965 138.235 88.135 ;
        RECT 138.525 87.965 138.695 88.135 ;
        RECT 138.985 87.965 139.155 88.135 ;
        RECT 50.665 85.245 50.835 85.415 ;
        RECT 51.125 85.245 51.295 85.415 ;
        RECT 51.585 85.245 51.755 85.415 ;
        RECT 52.045 85.245 52.215 85.415 ;
        RECT 52.505 85.245 52.675 85.415 ;
        RECT 52.965 85.245 53.135 85.415 ;
        RECT 53.425 85.245 53.595 85.415 ;
        RECT 53.885 85.245 54.055 85.415 ;
        RECT 54.345 85.245 54.515 85.415 ;
        RECT 54.805 85.245 54.975 85.415 ;
        RECT 55.265 85.245 55.435 85.415 ;
        RECT 55.725 85.245 55.895 85.415 ;
        RECT 56.185 85.245 56.355 85.415 ;
        RECT 56.645 85.245 56.815 85.415 ;
        RECT 57.105 85.245 57.275 85.415 ;
        RECT 57.565 85.245 57.735 85.415 ;
        RECT 58.025 85.245 58.195 85.415 ;
        RECT 58.485 85.245 58.655 85.415 ;
        RECT 58.945 85.245 59.115 85.415 ;
        RECT 59.405 85.245 59.575 85.415 ;
        RECT 59.865 85.245 60.035 85.415 ;
        RECT 60.325 85.245 60.495 85.415 ;
        RECT 60.785 85.245 60.955 85.415 ;
        RECT 61.245 85.245 61.415 85.415 ;
        RECT 61.705 85.245 61.875 85.415 ;
        RECT 62.165 85.245 62.335 85.415 ;
        RECT 62.625 85.245 62.795 85.415 ;
        RECT 63.085 85.245 63.255 85.415 ;
        RECT 63.545 85.245 63.715 85.415 ;
        RECT 64.005 85.245 64.175 85.415 ;
        RECT 64.465 85.245 64.635 85.415 ;
        RECT 64.925 85.245 65.095 85.415 ;
        RECT 65.385 85.245 65.555 85.415 ;
        RECT 65.845 85.245 66.015 85.415 ;
        RECT 66.305 85.245 66.475 85.415 ;
        RECT 66.765 85.245 66.935 85.415 ;
        RECT 67.225 85.245 67.395 85.415 ;
        RECT 67.685 85.245 67.855 85.415 ;
        RECT 68.145 85.245 68.315 85.415 ;
        RECT 68.605 85.245 68.775 85.415 ;
        RECT 69.065 85.245 69.235 85.415 ;
        RECT 69.525 85.245 69.695 85.415 ;
        RECT 69.985 85.245 70.155 85.415 ;
        RECT 70.445 85.245 70.615 85.415 ;
        RECT 70.905 85.245 71.075 85.415 ;
        RECT 71.365 85.245 71.535 85.415 ;
        RECT 71.825 85.245 71.995 85.415 ;
        RECT 72.285 85.245 72.455 85.415 ;
        RECT 72.745 85.245 72.915 85.415 ;
        RECT 73.205 85.245 73.375 85.415 ;
        RECT 73.665 85.245 73.835 85.415 ;
        RECT 74.125 85.245 74.295 85.415 ;
        RECT 74.585 85.245 74.755 85.415 ;
        RECT 75.045 85.245 75.215 85.415 ;
        RECT 75.505 85.245 75.675 85.415 ;
        RECT 75.965 85.245 76.135 85.415 ;
        RECT 76.425 85.245 76.595 85.415 ;
        RECT 76.885 85.245 77.055 85.415 ;
        RECT 77.345 85.245 77.515 85.415 ;
        RECT 77.805 85.245 77.975 85.415 ;
        RECT 78.265 85.245 78.435 85.415 ;
        RECT 78.725 85.245 78.895 85.415 ;
        RECT 79.185 85.245 79.355 85.415 ;
        RECT 79.645 85.245 79.815 85.415 ;
        RECT 80.105 85.245 80.275 85.415 ;
        RECT 80.565 85.245 80.735 85.415 ;
        RECT 81.025 85.245 81.195 85.415 ;
        RECT 81.485 85.245 81.655 85.415 ;
        RECT 81.945 85.245 82.115 85.415 ;
        RECT 82.405 85.245 82.575 85.415 ;
        RECT 82.865 85.245 83.035 85.415 ;
        RECT 83.325 85.245 83.495 85.415 ;
        RECT 83.785 85.245 83.955 85.415 ;
        RECT 84.245 85.245 84.415 85.415 ;
        RECT 84.705 85.245 84.875 85.415 ;
        RECT 85.165 85.245 85.335 85.415 ;
        RECT 85.625 85.245 85.795 85.415 ;
        RECT 86.085 85.245 86.255 85.415 ;
        RECT 86.545 85.245 86.715 85.415 ;
        RECT 87.005 85.245 87.175 85.415 ;
        RECT 87.465 85.245 87.635 85.415 ;
        RECT 87.925 85.245 88.095 85.415 ;
        RECT 88.385 85.245 88.555 85.415 ;
        RECT 88.845 85.245 89.015 85.415 ;
        RECT 89.305 85.245 89.475 85.415 ;
        RECT 89.765 85.245 89.935 85.415 ;
        RECT 90.225 85.245 90.395 85.415 ;
        RECT 90.685 85.245 90.855 85.415 ;
        RECT 91.145 85.245 91.315 85.415 ;
        RECT 91.605 85.245 91.775 85.415 ;
        RECT 92.065 85.245 92.235 85.415 ;
        RECT 92.525 85.245 92.695 85.415 ;
        RECT 92.985 85.245 93.155 85.415 ;
        RECT 93.445 85.245 93.615 85.415 ;
        RECT 93.905 85.245 94.075 85.415 ;
        RECT 94.365 85.245 94.535 85.415 ;
        RECT 94.825 85.245 94.995 85.415 ;
        RECT 95.285 85.245 95.455 85.415 ;
        RECT 95.745 85.245 95.915 85.415 ;
        RECT 96.205 85.245 96.375 85.415 ;
        RECT 96.665 85.245 96.835 85.415 ;
        RECT 97.125 85.245 97.295 85.415 ;
        RECT 97.585 85.245 97.755 85.415 ;
        RECT 98.045 85.245 98.215 85.415 ;
        RECT 98.505 85.245 98.675 85.415 ;
        RECT 98.965 85.245 99.135 85.415 ;
        RECT 99.425 85.245 99.595 85.415 ;
        RECT 99.885 85.245 100.055 85.415 ;
        RECT 100.345 85.245 100.515 85.415 ;
        RECT 100.805 85.245 100.975 85.415 ;
        RECT 101.265 85.245 101.435 85.415 ;
        RECT 101.725 85.245 101.895 85.415 ;
        RECT 102.185 85.245 102.355 85.415 ;
        RECT 102.645 85.245 102.815 85.415 ;
        RECT 103.105 85.245 103.275 85.415 ;
        RECT 103.565 85.245 103.735 85.415 ;
        RECT 104.025 85.245 104.195 85.415 ;
        RECT 104.485 85.245 104.655 85.415 ;
        RECT 104.945 85.245 105.115 85.415 ;
        RECT 105.405 85.245 105.575 85.415 ;
        RECT 105.865 85.245 106.035 85.415 ;
        RECT 106.325 85.245 106.495 85.415 ;
        RECT 106.785 85.245 106.955 85.415 ;
        RECT 107.245 85.245 107.415 85.415 ;
        RECT 107.705 85.245 107.875 85.415 ;
        RECT 108.165 85.245 108.335 85.415 ;
        RECT 108.625 85.245 108.795 85.415 ;
        RECT 109.085 85.245 109.255 85.415 ;
        RECT 109.545 85.245 109.715 85.415 ;
        RECT 110.005 85.245 110.175 85.415 ;
        RECT 110.465 85.245 110.635 85.415 ;
        RECT 110.925 85.245 111.095 85.415 ;
        RECT 111.385 85.245 111.555 85.415 ;
        RECT 111.845 85.245 112.015 85.415 ;
        RECT 112.305 85.245 112.475 85.415 ;
        RECT 112.765 85.245 112.935 85.415 ;
        RECT 113.225 85.245 113.395 85.415 ;
        RECT 113.685 85.245 113.855 85.415 ;
        RECT 114.145 85.245 114.315 85.415 ;
        RECT 114.605 85.245 114.775 85.415 ;
        RECT 115.065 85.245 115.235 85.415 ;
        RECT 115.525 85.245 115.695 85.415 ;
        RECT 115.985 85.245 116.155 85.415 ;
        RECT 116.445 85.245 116.615 85.415 ;
        RECT 116.905 85.245 117.075 85.415 ;
        RECT 117.365 85.245 117.535 85.415 ;
        RECT 117.825 85.245 117.995 85.415 ;
        RECT 118.285 85.245 118.455 85.415 ;
        RECT 118.745 85.245 118.915 85.415 ;
        RECT 119.205 85.245 119.375 85.415 ;
        RECT 119.665 85.245 119.835 85.415 ;
        RECT 120.125 85.245 120.295 85.415 ;
        RECT 120.585 85.245 120.755 85.415 ;
        RECT 121.045 85.245 121.215 85.415 ;
        RECT 121.505 85.245 121.675 85.415 ;
        RECT 121.965 85.245 122.135 85.415 ;
        RECT 122.425 85.245 122.595 85.415 ;
        RECT 122.885 85.245 123.055 85.415 ;
        RECT 123.345 85.245 123.515 85.415 ;
        RECT 123.805 85.245 123.975 85.415 ;
        RECT 124.265 85.245 124.435 85.415 ;
        RECT 124.725 85.245 124.895 85.415 ;
        RECT 125.185 85.245 125.355 85.415 ;
        RECT 125.645 85.245 125.815 85.415 ;
        RECT 126.105 85.245 126.275 85.415 ;
        RECT 126.565 85.245 126.735 85.415 ;
        RECT 127.025 85.245 127.195 85.415 ;
        RECT 127.485 85.245 127.655 85.415 ;
        RECT 127.945 85.245 128.115 85.415 ;
        RECT 128.405 85.245 128.575 85.415 ;
        RECT 128.865 85.245 129.035 85.415 ;
        RECT 129.325 85.245 129.495 85.415 ;
        RECT 129.785 85.245 129.955 85.415 ;
        RECT 130.245 85.245 130.415 85.415 ;
        RECT 130.705 85.245 130.875 85.415 ;
        RECT 131.165 85.245 131.335 85.415 ;
        RECT 131.625 85.245 131.795 85.415 ;
        RECT 132.085 85.245 132.255 85.415 ;
        RECT 132.545 85.245 132.715 85.415 ;
        RECT 133.005 85.245 133.175 85.415 ;
        RECT 133.465 85.245 133.635 85.415 ;
        RECT 133.925 85.245 134.095 85.415 ;
        RECT 134.385 85.245 134.555 85.415 ;
        RECT 134.845 85.245 135.015 85.415 ;
        RECT 135.305 85.245 135.475 85.415 ;
        RECT 135.765 85.245 135.935 85.415 ;
        RECT 136.225 85.245 136.395 85.415 ;
        RECT 136.685 85.245 136.855 85.415 ;
        RECT 137.145 85.245 137.315 85.415 ;
        RECT 137.605 85.245 137.775 85.415 ;
        RECT 138.065 85.245 138.235 85.415 ;
        RECT 138.525 85.245 138.695 85.415 ;
        RECT 138.985 85.245 139.155 85.415 ;
        RECT 50.665 82.525 50.835 82.695 ;
        RECT 51.125 82.525 51.295 82.695 ;
        RECT 51.585 82.525 51.755 82.695 ;
        RECT 52.045 82.525 52.215 82.695 ;
        RECT 52.505 82.525 52.675 82.695 ;
        RECT 52.965 82.525 53.135 82.695 ;
        RECT 53.425 82.525 53.595 82.695 ;
        RECT 53.885 82.525 54.055 82.695 ;
        RECT 54.345 82.525 54.515 82.695 ;
        RECT 54.805 82.525 54.975 82.695 ;
        RECT 55.265 82.525 55.435 82.695 ;
        RECT 55.725 82.525 55.895 82.695 ;
        RECT 56.185 82.525 56.355 82.695 ;
        RECT 56.645 82.525 56.815 82.695 ;
        RECT 57.105 82.525 57.275 82.695 ;
        RECT 57.565 82.525 57.735 82.695 ;
        RECT 58.025 82.525 58.195 82.695 ;
        RECT 58.485 82.525 58.655 82.695 ;
        RECT 58.945 82.525 59.115 82.695 ;
        RECT 59.405 82.525 59.575 82.695 ;
        RECT 59.865 82.525 60.035 82.695 ;
        RECT 60.325 82.525 60.495 82.695 ;
        RECT 60.785 82.525 60.955 82.695 ;
        RECT 61.245 82.525 61.415 82.695 ;
        RECT 61.705 82.525 61.875 82.695 ;
        RECT 62.165 82.525 62.335 82.695 ;
        RECT 62.625 82.525 62.795 82.695 ;
        RECT 63.085 82.525 63.255 82.695 ;
        RECT 63.545 82.525 63.715 82.695 ;
        RECT 64.005 82.525 64.175 82.695 ;
        RECT 64.465 82.525 64.635 82.695 ;
        RECT 64.925 82.525 65.095 82.695 ;
        RECT 65.385 82.525 65.555 82.695 ;
        RECT 65.845 82.525 66.015 82.695 ;
        RECT 66.305 82.525 66.475 82.695 ;
        RECT 66.765 82.525 66.935 82.695 ;
        RECT 67.225 82.525 67.395 82.695 ;
        RECT 67.685 82.525 67.855 82.695 ;
        RECT 68.145 82.525 68.315 82.695 ;
        RECT 68.605 82.525 68.775 82.695 ;
        RECT 69.065 82.525 69.235 82.695 ;
        RECT 69.525 82.525 69.695 82.695 ;
        RECT 69.985 82.525 70.155 82.695 ;
        RECT 70.445 82.525 70.615 82.695 ;
        RECT 70.905 82.525 71.075 82.695 ;
        RECT 71.365 82.525 71.535 82.695 ;
        RECT 71.825 82.525 71.995 82.695 ;
        RECT 72.285 82.525 72.455 82.695 ;
        RECT 72.745 82.525 72.915 82.695 ;
        RECT 73.205 82.525 73.375 82.695 ;
        RECT 73.665 82.525 73.835 82.695 ;
        RECT 74.125 82.525 74.295 82.695 ;
        RECT 74.585 82.525 74.755 82.695 ;
        RECT 75.045 82.525 75.215 82.695 ;
        RECT 75.505 82.525 75.675 82.695 ;
        RECT 75.965 82.525 76.135 82.695 ;
        RECT 76.425 82.525 76.595 82.695 ;
        RECT 76.885 82.525 77.055 82.695 ;
        RECT 77.345 82.525 77.515 82.695 ;
        RECT 77.805 82.525 77.975 82.695 ;
        RECT 78.265 82.525 78.435 82.695 ;
        RECT 78.725 82.525 78.895 82.695 ;
        RECT 79.185 82.525 79.355 82.695 ;
        RECT 79.645 82.525 79.815 82.695 ;
        RECT 80.105 82.525 80.275 82.695 ;
        RECT 80.565 82.525 80.735 82.695 ;
        RECT 81.025 82.525 81.195 82.695 ;
        RECT 81.485 82.525 81.655 82.695 ;
        RECT 81.945 82.525 82.115 82.695 ;
        RECT 82.405 82.525 82.575 82.695 ;
        RECT 82.865 82.525 83.035 82.695 ;
        RECT 83.325 82.525 83.495 82.695 ;
        RECT 83.785 82.525 83.955 82.695 ;
        RECT 84.245 82.525 84.415 82.695 ;
        RECT 84.705 82.525 84.875 82.695 ;
        RECT 85.165 82.525 85.335 82.695 ;
        RECT 85.625 82.525 85.795 82.695 ;
        RECT 86.085 82.525 86.255 82.695 ;
        RECT 86.545 82.525 86.715 82.695 ;
        RECT 87.005 82.525 87.175 82.695 ;
        RECT 87.465 82.525 87.635 82.695 ;
        RECT 87.925 82.525 88.095 82.695 ;
        RECT 88.385 82.525 88.555 82.695 ;
        RECT 88.845 82.525 89.015 82.695 ;
        RECT 89.305 82.525 89.475 82.695 ;
        RECT 89.765 82.525 89.935 82.695 ;
        RECT 90.225 82.525 90.395 82.695 ;
        RECT 90.685 82.525 90.855 82.695 ;
        RECT 91.145 82.525 91.315 82.695 ;
        RECT 91.605 82.525 91.775 82.695 ;
        RECT 92.065 82.525 92.235 82.695 ;
        RECT 92.525 82.525 92.695 82.695 ;
        RECT 92.985 82.525 93.155 82.695 ;
        RECT 93.445 82.525 93.615 82.695 ;
        RECT 93.905 82.525 94.075 82.695 ;
        RECT 94.365 82.525 94.535 82.695 ;
        RECT 94.825 82.525 94.995 82.695 ;
        RECT 95.285 82.525 95.455 82.695 ;
        RECT 95.745 82.525 95.915 82.695 ;
        RECT 96.205 82.525 96.375 82.695 ;
        RECT 96.665 82.525 96.835 82.695 ;
        RECT 97.125 82.525 97.295 82.695 ;
        RECT 97.585 82.525 97.755 82.695 ;
        RECT 98.045 82.525 98.215 82.695 ;
        RECT 98.505 82.525 98.675 82.695 ;
        RECT 98.965 82.525 99.135 82.695 ;
        RECT 99.425 82.525 99.595 82.695 ;
        RECT 99.885 82.525 100.055 82.695 ;
        RECT 100.345 82.525 100.515 82.695 ;
        RECT 100.805 82.525 100.975 82.695 ;
        RECT 101.265 82.525 101.435 82.695 ;
        RECT 101.725 82.525 101.895 82.695 ;
        RECT 102.185 82.525 102.355 82.695 ;
        RECT 102.645 82.525 102.815 82.695 ;
        RECT 103.105 82.525 103.275 82.695 ;
        RECT 103.565 82.525 103.735 82.695 ;
        RECT 104.025 82.525 104.195 82.695 ;
        RECT 104.485 82.525 104.655 82.695 ;
        RECT 104.945 82.525 105.115 82.695 ;
        RECT 105.405 82.525 105.575 82.695 ;
        RECT 105.865 82.525 106.035 82.695 ;
        RECT 106.325 82.525 106.495 82.695 ;
        RECT 106.785 82.525 106.955 82.695 ;
        RECT 107.245 82.525 107.415 82.695 ;
        RECT 107.705 82.525 107.875 82.695 ;
        RECT 108.165 82.525 108.335 82.695 ;
        RECT 108.625 82.525 108.795 82.695 ;
        RECT 109.085 82.525 109.255 82.695 ;
        RECT 109.545 82.525 109.715 82.695 ;
        RECT 110.005 82.525 110.175 82.695 ;
        RECT 110.465 82.525 110.635 82.695 ;
        RECT 110.925 82.525 111.095 82.695 ;
        RECT 111.385 82.525 111.555 82.695 ;
        RECT 111.845 82.525 112.015 82.695 ;
        RECT 112.305 82.525 112.475 82.695 ;
        RECT 112.765 82.525 112.935 82.695 ;
        RECT 113.225 82.525 113.395 82.695 ;
        RECT 113.685 82.525 113.855 82.695 ;
        RECT 114.145 82.525 114.315 82.695 ;
        RECT 114.605 82.525 114.775 82.695 ;
        RECT 115.065 82.525 115.235 82.695 ;
        RECT 115.525 82.525 115.695 82.695 ;
        RECT 115.985 82.525 116.155 82.695 ;
        RECT 116.445 82.525 116.615 82.695 ;
        RECT 116.905 82.525 117.075 82.695 ;
        RECT 117.365 82.525 117.535 82.695 ;
        RECT 117.825 82.525 117.995 82.695 ;
        RECT 118.285 82.525 118.455 82.695 ;
        RECT 118.745 82.525 118.915 82.695 ;
        RECT 119.205 82.525 119.375 82.695 ;
        RECT 119.665 82.525 119.835 82.695 ;
        RECT 120.125 82.525 120.295 82.695 ;
        RECT 120.585 82.525 120.755 82.695 ;
        RECT 121.045 82.525 121.215 82.695 ;
        RECT 121.505 82.525 121.675 82.695 ;
        RECT 121.965 82.525 122.135 82.695 ;
        RECT 122.425 82.525 122.595 82.695 ;
        RECT 122.885 82.525 123.055 82.695 ;
        RECT 123.345 82.525 123.515 82.695 ;
        RECT 123.805 82.525 123.975 82.695 ;
        RECT 124.265 82.525 124.435 82.695 ;
        RECT 124.725 82.525 124.895 82.695 ;
        RECT 125.185 82.525 125.355 82.695 ;
        RECT 125.645 82.525 125.815 82.695 ;
        RECT 126.105 82.525 126.275 82.695 ;
        RECT 126.565 82.525 126.735 82.695 ;
        RECT 127.025 82.525 127.195 82.695 ;
        RECT 127.485 82.525 127.655 82.695 ;
        RECT 127.945 82.525 128.115 82.695 ;
        RECT 128.405 82.525 128.575 82.695 ;
        RECT 128.865 82.525 129.035 82.695 ;
        RECT 129.325 82.525 129.495 82.695 ;
        RECT 129.785 82.525 129.955 82.695 ;
        RECT 130.245 82.525 130.415 82.695 ;
        RECT 130.705 82.525 130.875 82.695 ;
        RECT 131.165 82.525 131.335 82.695 ;
        RECT 131.625 82.525 131.795 82.695 ;
        RECT 132.085 82.525 132.255 82.695 ;
        RECT 132.545 82.525 132.715 82.695 ;
        RECT 133.005 82.525 133.175 82.695 ;
        RECT 133.465 82.525 133.635 82.695 ;
        RECT 133.925 82.525 134.095 82.695 ;
        RECT 134.385 82.525 134.555 82.695 ;
        RECT 134.845 82.525 135.015 82.695 ;
        RECT 135.305 82.525 135.475 82.695 ;
        RECT 135.765 82.525 135.935 82.695 ;
        RECT 136.225 82.525 136.395 82.695 ;
        RECT 136.685 82.525 136.855 82.695 ;
        RECT 137.145 82.525 137.315 82.695 ;
        RECT 137.605 82.525 137.775 82.695 ;
        RECT 138.065 82.525 138.235 82.695 ;
        RECT 138.525 82.525 138.695 82.695 ;
        RECT 138.985 82.525 139.155 82.695 ;
        RECT 50.665 79.805 50.835 79.975 ;
        RECT 51.125 79.805 51.295 79.975 ;
        RECT 51.585 79.805 51.755 79.975 ;
        RECT 52.045 79.805 52.215 79.975 ;
        RECT 52.505 79.805 52.675 79.975 ;
        RECT 52.965 79.805 53.135 79.975 ;
        RECT 53.425 79.805 53.595 79.975 ;
        RECT 53.885 79.805 54.055 79.975 ;
        RECT 54.345 79.805 54.515 79.975 ;
        RECT 54.805 79.805 54.975 79.975 ;
        RECT 55.265 79.805 55.435 79.975 ;
        RECT 55.725 79.805 55.895 79.975 ;
        RECT 56.185 79.805 56.355 79.975 ;
        RECT 56.645 79.805 56.815 79.975 ;
        RECT 57.105 79.805 57.275 79.975 ;
        RECT 57.565 79.805 57.735 79.975 ;
        RECT 58.025 79.805 58.195 79.975 ;
        RECT 58.485 79.805 58.655 79.975 ;
        RECT 58.945 79.805 59.115 79.975 ;
        RECT 59.405 79.805 59.575 79.975 ;
        RECT 59.865 79.805 60.035 79.975 ;
        RECT 60.325 79.805 60.495 79.975 ;
        RECT 60.785 79.805 60.955 79.975 ;
        RECT 61.245 79.805 61.415 79.975 ;
        RECT 61.705 79.805 61.875 79.975 ;
        RECT 62.165 79.805 62.335 79.975 ;
        RECT 62.625 79.805 62.795 79.975 ;
        RECT 63.085 79.805 63.255 79.975 ;
        RECT 63.545 79.805 63.715 79.975 ;
        RECT 64.005 79.805 64.175 79.975 ;
        RECT 64.465 79.805 64.635 79.975 ;
        RECT 64.925 79.805 65.095 79.975 ;
        RECT 65.385 79.805 65.555 79.975 ;
        RECT 65.845 79.805 66.015 79.975 ;
        RECT 66.305 79.805 66.475 79.975 ;
        RECT 66.765 79.805 66.935 79.975 ;
        RECT 67.225 79.805 67.395 79.975 ;
        RECT 67.685 79.805 67.855 79.975 ;
        RECT 68.145 79.805 68.315 79.975 ;
        RECT 68.605 79.805 68.775 79.975 ;
        RECT 69.065 79.805 69.235 79.975 ;
        RECT 69.525 79.805 69.695 79.975 ;
        RECT 69.985 79.805 70.155 79.975 ;
        RECT 70.445 79.805 70.615 79.975 ;
        RECT 70.905 79.805 71.075 79.975 ;
        RECT 71.365 79.805 71.535 79.975 ;
        RECT 71.825 79.805 71.995 79.975 ;
        RECT 72.285 79.805 72.455 79.975 ;
        RECT 72.745 79.805 72.915 79.975 ;
        RECT 73.205 79.805 73.375 79.975 ;
        RECT 73.665 79.805 73.835 79.975 ;
        RECT 74.125 79.805 74.295 79.975 ;
        RECT 74.585 79.805 74.755 79.975 ;
        RECT 75.045 79.805 75.215 79.975 ;
        RECT 75.505 79.805 75.675 79.975 ;
        RECT 75.965 79.805 76.135 79.975 ;
        RECT 76.425 79.805 76.595 79.975 ;
        RECT 76.885 79.805 77.055 79.975 ;
        RECT 77.345 79.805 77.515 79.975 ;
        RECT 77.805 79.805 77.975 79.975 ;
        RECT 78.265 79.805 78.435 79.975 ;
        RECT 78.725 79.805 78.895 79.975 ;
        RECT 79.185 79.805 79.355 79.975 ;
        RECT 79.645 79.805 79.815 79.975 ;
        RECT 80.105 79.805 80.275 79.975 ;
        RECT 80.565 79.805 80.735 79.975 ;
        RECT 81.025 79.805 81.195 79.975 ;
        RECT 81.485 79.805 81.655 79.975 ;
        RECT 81.945 79.805 82.115 79.975 ;
        RECT 82.405 79.805 82.575 79.975 ;
        RECT 82.865 79.805 83.035 79.975 ;
        RECT 83.325 79.805 83.495 79.975 ;
        RECT 83.785 79.805 83.955 79.975 ;
        RECT 84.245 79.805 84.415 79.975 ;
        RECT 84.705 79.805 84.875 79.975 ;
        RECT 85.165 79.805 85.335 79.975 ;
        RECT 85.625 79.805 85.795 79.975 ;
        RECT 86.085 79.805 86.255 79.975 ;
        RECT 86.545 79.805 86.715 79.975 ;
        RECT 87.005 79.805 87.175 79.975 ;
        RECT 87.465 79.805 87.635 79.975 ;
        RECT 87.925 79.805 88.095 79.975 ;
        RECT 88.385 79.805 88.555 79.975 ;
        RECT 88.845 79.805 89.015 79.975 ;
        RECT 89.305 79.805 89.475 79.975 ;
        RECT 89.765 79.805 89.935 79.975 ;
        RECT 90.225 79.805 90.395 79.975 ;
        RECT 90.685 79.805 90.855 79.975 ;
        RECT 91.145 79.805 91.315 79.975 ;
        RECT 91.605 79.805 91.775 79.975 ;
        RECT 92.065 79.805 92.235 79.975 ;
        RECT 92.525 79.805 92.695 79.975 ;
        RECT 92.985 79.805 93.155 79.975 ;
        RECT 93.445 79.805 93.615 79.975 ;
        RECT 93.905 79.805 94.075 79.975 ;
        RECT 94.365 79.805 94.535 79.975 ;
        RECT 94.825 79.805 94.995 79.975 ;
        RECT 95.285 79.805 95.455 79.975 ;
        RECT 95.745 79.805 95.915 79.975 ;
        RECT 96.205 79.805 96.375 79.975 ;
        RECT 96.665 79.805 96.835 79.975 ;
        RECT 97.125 79.805 97.295 79.975 ;
        RECT 97.585 79.805 97.755 79.975 ;
        RECT 98.045 79.805 98.215 79.975 ;
        RECT 98.505 79.805 98.675 79.975 ;
        RECT 98.965 79.805 99.135 79.975 ;
        RECT 99.425 79.805 99.595 79.975 ;
        RECT 99.885 79.805 100.055 79.975 ;
        RECT 100.345 79.805 100.515 79.975 ;
        RECT 100.805 79.805 100.975 79.975 ;
        RECT 101.265 79.805 101.435 79.975 ;
        RECT 101.725 79.805 101.895 79.975 ;
        RECT 102.185 79.805 102.355 79.975 ;
        RECT 102.645 79.805 102.815 79.975 ;
        RECT 103.105 79.805 103.275 79.975 ;
        RECT 103.565 79.805 103.735 79.975 ;
        RECT 104.025 79.805 104.195 79.975 ;
        RECT 104.485 79.805 104.655 79.975 ;
        RECT 104.945 79.805 105.115 79.975 ;
        RECT 105.405 79.805 105.575 79.975 ;
        RECT 105.865 79.805 106.035 79.975 ;
        RECT 106.325 79.805 106.495 79.975 ;
        RECT 106.785 79.805 106.955 79.975 ;
        RECT 107.245 79.805 107.415 79.975 ;
        RECT 107.705 79.805 107.875 79.975 ;
        RECT 108.165 79.805 108.335 79.975 ;
        RECT 108.625 79.805 108.795 79.975 ;
        RECT 109.085 79.805 109.255 79.975 ;
        RECT 109.545 79.805 109.715 79.975 ;
        RECT 110.005 79.805 110.175 79.975 ;
        RECT 110.465 79.805 110.635 79.975 ;
        RECT 110.925 79.805 111.095 79.975 ;
        RECT 111.385 79.805 111.555 79.975 ;
        RECT 111.845 79.805 112.015 79.975 ;
        RECT 112.305 79.805 112.475 79.975 ;
        RECT 112.765 79.805 112.935 79.975 ;
        RECT 113.225 79.805 113.395 79.975 ;
        RECT 113.685 79.805 113.855 79.975 ;
        RECT 114.145 79.805 114.315 79.975 ;
        RECT 114.605 79.805 114.775 79.975 ;
        RECT 115.065 79.805 115.235 79.975 ;
        RECT 115.525 79.805 115.695 79.975 ;
        RECT 115.985 79.805 116.155 79.975 ;
        RECT 116.445 79.805 116.615 79.975 ;
        RECT 116.905 79.805 117.075 79.975 ;
        RECT 117.365 79.805 117.535 79.975 ;
        RECT 117.825 79.805 117.995 79.975 ;
        RECT 118.285 79.805 118.455 79.975 ;
        RECT 118.745 79.805 118.915 79.975 ;
        RECT 119.205 79.805 119.375 79.975 ;
        RECT 119.665 79.805 119.835 79.975 ;
        RECT 120.125 79.805 120.295 79.975 ;
        RECT 120.585 79.805 120.755 79.975 ;
        RECT 121.045 79.805 121.215 79.975 ;
        RECT 121.505 79.805 121.675 79.975 ;
        RECT 121.965 79.805 122.135 79.975 ;
        RECT 122.425 79.805 122.595 79.975 ;
        RECT 122.885 79.805 123.055 79.975 ;
        RECT 123.345 79.805 123.515 79.975 ;
        RECT 123.805 79.805 123.975 79.975 ;
        RECT 124.265 79.805 124.435 79.975 ;
        RECT 124.725 79.805 124.895 79.975 ;
        RECT 125.185 79.805 125.355 79.975 ;
        RECT 125.645 79.805 125.815 79.975 ;
        RECT 126.105 79.805 126.275 79.975 ;
        RECT 126.565 79.805 126.735 79.975 ;
        RECT 127.025 79.805 127.195 79.975 ;
        RECT 127.485 79.805 127.655 79.975 ;
        RECT 127.945 79.805 128.115 79.975 ;
        RECT 128.405 79.805 128.575 79.975 ;
        RECT 128.865 79.805 129.035 79.975 ;
        RECT 129.325 79.805 129.495 79.975 ;
        RECT 129.785 79.805 129.955 79.975 ;
        RECT 130.245 79.805 130.415 79.975 ;
        RECT 130.705 79.805 130.875 79.975 ;
        RECT 131.165 79.805 131.335 79.975 ;
        RECT 131.625 79.805 131.795 79.975 ;
        RECT 132.085 79.805 132.255 79.975 ;
        RECT 132.545 79.805 132.715 79.975 ;
        RECT 133.005 79.805 133.175 79.975 ;
        RECT 133.465 79.805 133.635 79.975 ;
        RECT 133.925 79.805 134.095 79.975 ;
        RECT 134.385 79.805 134.555 79.975 ;
        RECT 134.845 79.805 135.015 79.975 ;
        RECT 135.305 79.805 135.475 79.975 ;
        RECT 135.765 79.805 135.935 79.975 ;
        RECT 136.225 79.805 136.395 79.975 ;
        RECT 136.685 79.805 136.855 79.975 ;
        RECT 137.145 79.805 137.315 79.975 ;
        RECT 137.605 79.805 137.775 79.975 ;
        RECT 138.065 79.805 138.235 79.975 ;
        RECT 138.525 79.805 138.695 79.975 ;
        RECT 138.985 79.805 139.155 79.975 ;
        RECT 50.665 77.085 50.835 77.255 ;
        RECT 51.125 77.085 51.295 77.255 ;
        RECT 51.585 77.085 51.755 77.255 ;
        RECT 52.045 77.085 52.215 77.255 ;
        RECT 52.505 77.085 52.675 77.255 ;
        RECT 52.965 77.085 53.135 77.255 ;
        RECT 53.425 77.085 53.595 77.255 ;
        RECT 53.885 77.085 54.055 77.255 ;
        RECT 54.345 77.085 54.515 77.255 ;
        RECT 54.805 77.085 54.975 77.255 ;
        RECT 55.265 77.085 55.435 77.255 ;
        RECT 55.725 77.085 55.895 77.255 ;
        RECT 56.185 77.085 56.355 77.255 ;
        RECT 56.645 77.085 56.815 77.255 ;
        RECT 57.105 77.085 57.275 77.255 ;
        RECT 57.565 77.085 57.735 77.255 ;
        RECT 58.025 77.085 58.195 77.255 ;
        RECT 58.485 77.085 58.655 77.255 ;
        RECT 58.945 77.085 59.115 77.255 ;
        RECT 59.405 77.085 59.575 77.255 ;
        RECT 59.865 77.085 60.035 77.255 ;
        RECT 60.325 77.085 60.495 77.255 ;
        RECT 60.785 77.085 60.955 77.255 ;
        RECT 61.245 77.085 61.415 77.255 ;
        RECT 61.705 77.085 61.875 77.255 ;
        RECT 62.165 77.085 62.335 77.255 ;
        RECT 62.625 77.085 62.795 77.255 ;
        RECT 63.085 77.085 63.255 77.255 ;
        RECT 63.545 77.085 63.715 77.255 ;
        RECT 64.005 77.085 64.175 77.255 ;
        RECT 64.465 77.085 64.635 77.255 ;
        RECT 64.925 77.085 65.095 77.255 ;
        RECT 65.385 77.085 65.555 77.255 ;
        RECT 65.845 77.085 66.015 77.255 ;
        RECT 66.305 77.085 66.475 77.255 ;
        RECT 66.765 77.085 66.935 77.255 ;
        RECT 67.225 77.085 67.395 77.255 ;
        RECT 67.685 77.085 67.855 77.255 ;
        RECT 68.145 77.085 68.315 77.255 ;
        RECT 68.605 77.085 68.775 77.255 ;
        RECT 69.065 77.085 69.235 77.255 ;
        RECT 69.525 77.085 69.695 77.255 ;
        RECT 69.985 77.085 70.155 77.255 ;
        RECT 70.445 77.085 70.615 77.255 ;
        RECT 70.905 77.085 71.075 77.255 ;
        RECT 71.365 77.085 71.535 77.255 ;
        RECT 71.825 77.085 71.995 77.255 ;
        RECT 72.285 77.085 72.455 77.255 ;
        RECT 72.745 77.085 72.915 77.255 ;
        RECT 73.205 77.085 73.375 77.255 ;
        RECT 73.665 77.085 73.835 77.255 ;
        RECT 74.125 77.085 74.295 77.255 ;
        RECT 74.585 77.085 74.755 77.255 ;
        RECT 75.045 77.085 75.215 77.255 ;
        RECT 75.505 77.085 75.675 77.255 ;
        RECT 75.965 77.085 76.135 77.255 ;
        RECT 76.425 77.085 76.595 77.255 ;
        RECT 76.885 77.085 77.055 77.255 ;
        RECT 77.345 77.085 77.515 77.255 ;
        RECT 77.805 77.085 77.975 77.255 ;
        RECT 78.265 77.085 78.435 77.255 ;
        RECT 78.725 77.085 78.895 77.255 ;
        RECT 79.185 77.085 79.355 77.255 ;
        RECT 79.645 77.085 79.815 77.255 ;
        RECT 80.105 77.085 80.275 77.255 ;
        RECT 80.565 77.085 80.735 77.255 ;
        RECT 81.025 77.085 81.195 77.255 ;
        RECT 81.485 77.085 81.655 77.255 ;
        RECT 81.945 77.085 82.115 77.255 ;
        RECT 82.405 77.085 82.575 77.255 ;
        RECT 82.865 77.085 83.035 77.255 ;
        RECT 83.325 77.085 83.495 77.255 ;
        RECT 83.785 77.085 83.955 77.255 ;
        RECT 84.245 77.085 84.415 77.255 ;
        RECT 84.705 77.085 84.875 77.255 ;
        RECT 85.165 77.085 85.335 77.255 ;
        RECT 85.625 77.085 85.795 77.255 ;
        RECT 86.085 77.085 86.255 77.255 ;
        RECT 86.545 77.085 86.715 77.255 ;
        RECT 87.005 77.085 87.175 77.255 ;
        RECT 87.465 77.085 87.635 77.255 ;
        RECT 87.925 77.085 88.095 77.255 ;
        RECT 88.385 77.085 88.555 77.255 ;
        RECT 88.845 77.085 89.015 77.255 ;
        RECT 89.305 77.085 89.475 77.255 ;
        RECT 89.765 77.085 89.935 77.255 ;
        RECT 90.225 77.085 90.395 77.255 ;
        RECT 90.685 77.085 90.855 77.255 ;
        RECT 91.145 77.085 91.315 77.255 ;
        RECT 91.605 77.085 91.775 77.255 ;
        RECT 92.065 77.085 92.235 77.255 ;
        RECT 92.525 77.085 92.695 77.255 ;
        RECT 92.985 77.085 93.155 77.255 ;
        RECT 93.445 77.085 93.615 77.255 ;
        RECT 93.905 77.085 94.075 77.255 ;
        RECT 94.365 77.085 94.535 77.255 ;
        RECT 94.825 77.085 94.995 77.255 ;
        RECT 95.285 77.085 95.455 77.255 ;
        RECT 95.745 77.085 95.915 77.255 ;
        RECT 96.205 77.085 96.375 77.255 ;
        RECT 96.665 77.085 96.835 77.255 ;
        RECT 97.125 77.085 97.295 77.255 ;
        RECT 97.585 77.085 97.755 77.255 ;
        RECT 98.045 77.085 98.215 77.255 ;
        RECT 98.505 77.085 98.675 77.255 ;
        RECT 98.965 77.085 99.135 77.255 ;
        RECT 99.425 77.085 99.595 77.255 ;
        RECT 99.885 77.085 100.055 77.255 ;
        RECT 100.345 77.085 100.515 77.255 ;
        RECT 100.805 77.085 100.975 77.255 ;
        RECT 101.265 77.085 101.435 77.255 ;
        RECT 101.725 77.085 101.895 77.255 ;
        RECT 102.185 77.085 102.355 77.255 ;
        RECT 102.645 77.085 102.815 77.255 ;
        RECT 103.105 77.085 103.275 77.255 ;
        RECT 103.565 77.085 103.735 77.255 ;
        RECT 104.025 77.085 104.195 77.255 ;
        RECT 104.485 77.085 104.655 77.255 ;
        RECT 104.945 77.085 105.115 77.255 ;
        RECT 105.405 77.085 105.575 77.255 ;
        RECT 105.865 77.085 106.035 77.255 ;
        RECT 106.325 77.085 106.495 77.255 ;
        RECT 106.785 77.085 106.955 77.255 ;
        RECT 107.245 77.085 107.415 77.255 ;
        RECT 107.705 77.085 107.875 77.255 ;
        RECT 108.165 77.085 108.335 77.255 ;
        RECT 108.625 77.085 108.795 77.255 ;
        RECT 109.085 77.085 109.255 77.255 ;
        RECT 109.545 77.085 109.715 77.255 ;
        RECT 110.005 77.085 110.175 77.255 ;
        RECT 110.465 77.085 110.635 77.255 ;
        RECT 110.925 77.085 111.095 77.255 ;
        RECT 111.385 77.085 111.555 77.255 ;
        RECT 111.845 77.085 112.015 77.255 ;
        RECT 112.305 77.085 112.475 77.255 ;
        RECT 112.765 77.085 112.935 77.255 ;
        RECT 113.225 77.085 113.395 77.255 ;
        RECT 113.685 77.085 113.855 77.255 ;
        RECT 114.145 77.085 114.315 77.255 ;
        RECT 114.605 77.085 114.775 77.255 ;
        RECT 115.065 77.085 115.235 77.255 ;
        RECT 115.525 77.085 115.695 77.255 ;
        RECT 115.985 77.085 116.155 77.255 ;
        RECT 116.445 77.085 116.615 77.255 ;
        RECT 116.905 77.085 117.075 77.255 ;
        RECT 117.365 77.085 117.535 77.255 ;
        RECT 117.825 77.085 117.995 77.255 ;
        RECT 118.285 77.085 118.455 77.255 ;
        RECT 118.745 77.085 118.915 77.255 ;
        RECT 119.205 77.085 119.375 77.255 ;
        RECT 119.665 77.085 119.835 77.255 ;
        RECT 120.125 77.085 120.295 77.255 ;
        RECT 120.585 77.085 120.755 77.255 ;
        RECT 121.045 77.085 121.215 77.255 ;
        RECT 121.505 77.085 121.675 77.255 ;
        RECT 121.965 77.085 122.135 77.255 ;
        RECT 122.425 77.085 122.595 77.255 ;
        RECT 122.885 77.085 123.055 77.255 ;
        RECT 123.345 77.085 123.515 77.255 ;
        RECT 123.805 77.085 123.975 77.255 ;
        RECT 124.265 77.085 124.435 77.255 ;
        RECT 124.725 77.085 124.895 77.255 ;
        RECT 125.185 77.085 125.355 77.255 ;
        RECT 125.645 77.085 125.815 77.255 ;
        RECT 126.105 77.085 126.275 77.255 ;
        RECT 126.565 77.085 126.735 77.255 ;
        RECT 127.025 77.085 127.195 77.255 ;
        RECT 127.485 77.085 127.655 77.255 ;
        RECT 127.945 77.085 128.115 77.255 ;
        RECT 128.405 77.085 128.575 77.255 ;
        RECT 128.865 77.085 129.035 77.255 ;
        RECT 129.325 77.085 129.495 77.255 ;
        RECT 129.785 77.085 129.955 77.255 ;
        RECT 130.245 77.085 130.415 77.255 ;
        RECT 130.705 77.085 130.875 77.255 ;
        RECT 131.165 77.085 131.335 77.255 ;
        RECT 131.625 77.085 131.795 77.255 ;
        RECT 132.085 77.085 132.255 77.255 ;
        RECT 132.545 77.085 132.715 77.255 ;
        RECT 133.005 77.085 133.175 77.255 ;
        RECT 133.465 77.085 133.635 77.255 ;
        RECT 133.925 77.085 134.095 77.255 ;
        RECT 134.385 77.085 134.555 77.255 ;
        RECT 134.845 77.085 135.015 77.255 ;
        RECT 135.305 77.085 135.475 77.255 ;
        RECT 135.765 77.085 135.935 77.255 ;
        RECT 136.225 77.085 136.395 77.255 ;
        RECT 136.685 77.085 136.855 77.255 ;
        RECT 137.145 77.085 137.315 77.255 ;
        RECT 137.605 77.085 137.775 77.255 ;
        RECT 138.065 77.085 138.235 77.255 ;
        RECT 138.525 77.085 138.695 77.255 ;
        RECT 138.985 77.085 139.155 77.255 ;
        RECT 50.665 74.365 50.835 74.535 ;
        RECT 51.125 74.365 51.295 74.535 ;
        RECT 51.585 74.365 51.755 74.535 ;
        RECT 52.045 74.365 52.215 74.535 ;
        RECT 52.505 74.365 52.675 74.535 ;
        RECT 52.965 74.365 53.135 74.535 ;
        RECT 53.425 74.365 53.595 74.535 ;
        RECT 53.885 74.365 54.055 74.535 ;
        RECT 54.345 74.365 54.515 74.535 ;
        RECT 54.805 74.365 54.975 74.535 ;
        RECT 55.265 74.365 55.435 74.535 ;
        RECT 55.725 74.365 55.895 74.535 ;
        RECT 56.185 74.365 56.355 74.535 ;
        RECT 56.645 74.365 56.815 74.535 ;
        RECT 57.105 74.365 57.275 74.535 ;
        RECT 57.565 74.365 57.735 74.535 ;
        RECT 58.025 74.365 58.195 74.535 ;
        RECT 58.485 74.365 58.655 74.535 ;
        RECT 58.945 74.365 59.115 74.535 ;
        RECT 59.405 74.365 59.575 74.535 ;
        RECT 59.865 74.365 60.035 74.535 ;
        RECT 60.325 74.365 60.495 74.535 ;
        RECT 60.785 74.365 60.955 74.535 ;
        RECT 61.245 74.365 61.415 74.535 ;
        RECT 61.705 74.365 61.875 74.535 ;
        RECT 62.165 74.365 62.335 74.535 ;
        RECT 62.625 74.365 62.795 74.535 ;
        RECT 63.085 74.365 63.255 74.535 ;
        RECT 63.545 74.365 63.715 74.535 ;
        RECT 64.005 74.365 64.175 74.535 ;
        RECT 64.465 74.365 64.635 74.535 ;
        RECT 64.925 74.365 65.095 74.535 ;
        RECT 65.385 74.365 65.555 74.535 ;
        RECT 65.845 74.365 66.015 74.535 ;
        RECT 66.305 74.365 66.475 74.535 ;
        RECT 66.765 74.365 66.935 74.535 ;
        RECT 67.225 74.365 67.395 74.535 ;
        RECT 67.685 74.365 67.855 74.535 ;
        RECT 68.145 74.365 68.315 74.535 ;
        RECT 68.605 74.365 68.775 74.535 ;
        RECT 69.065 74.365 69.235 74.535 ;
        RECT 69.525 74.365 69.695 74.535 ;
        RECT 69.985 74.365 70.155 74.535 ;
        RECT 70.445 74.365 70.615 74.535 ;
        RECT 70.905 74.365 71.075 74.535 ;
        RECT 71.365 74.365 71.535 74.535 ;
        RECT 71.825 74.365 71.995 74.535 ;
        RECT 72.285 74.365 72.455 74.535 ;
        RECT 72.745 74.365 72.915 74.535 ;
        RECT 73.205 74.365 73.375 74.535 ;
        RECT 73.665 74.365 73.835 74.535 ;
        RECT 74.125 74.365 74.295 74.535 ;
        RECT 74.585 74.365 74.755 74.535 ;
        RECT 75.045 74.365 75.215 74.535 ;
        RECT 75.505 74.365 75.675 74.535 ;
        RECT 75.965 74.365 76.135 74.535 ;
        RECT 76.425 74.365 76.595 74.535 ;
        RECT 76.885 74.365 77.055 74.535 ;
        RECT 77.345 74.365 77.515 74.535 ;
        RECT 77.805 74.365 77.975 74.535 ;
        RECT 78.265 74.365 78.435 74.535 ;
        RECT 78.725 74.365 78.895 74.535 ;
        RECT 79.185 74.365 79.355 74.535 ;
        RECT 79.645 74.365 79.815 74.535 ;
        RECT 80.105 74.365 80.275 74.535 ;
        RECT 80.565 74.365 80.735 74.535 ;
        RECT 81.025 74.365 81.195 74.535 ;
        RECT 81.485 74.365 81.655 74.535 ;
        RECT 81.945 74.365 82.115 74.535 ;
        RECT 82.405 74.365 82.575 74.535 ;
        RECT 82.865 74.365 83.035 74.535 ;
        RECT 83.325 74.365 83.495 74.535 ;
        RECT 83.785 74.365 83.955 74.535 ;
        RECT 84.245 74.365 84.415 74.535 ;
        RECT 84.705 74.365 84.875 74.535 ;
        RECT 85.165 74.365 85.335 74.535 ;
        RECT 85.625 74.365 85.795 74.535 ;
        RECT 86.085 74.365 86.255 74.535 ;
        RECT 86.545 74.365 86.715 74.535 ;
        RECT 87.005 74.365 87.175 74.535 ;
        RECT 87.465 74.365 87.635 74.535 ;
        RECT 87.925 74.365 88.095 74.535 ;
        RECT 88.385 74.365 88.555 74.535 ;
        RECT 88.845 74.365 89.015 74.535 ;
        RECT 89.305 74.365 89.475 74.535 ;
        RECT 89.765 74.365 89.935 74.535 ;
        RECT 90.225 74.365 90.395 74.535 ;
        RECT 90.685 74.365 90.855 74.535 ;
        RECT 91.145 74.365 91.315 74.535 ;
        RECT 91.605 74.365 91.775 74.535 ;
        RECT 92.065 74.365 92.235 74.535 ;
        RECT 92.525 74.365 92.695 74.535 ;
        RECT 92.985 74.365 93.155 74.535 ;
        RECT 93.445 74.365 93.615 74.535 ;
        RECT 93.905 74.365 94.075 74.535 ;
        RECT 94.365 74.365 94.535 74.535 ;
        RECT 94.825 74.365 94.995 74.535 ;
        RECT 95.285 74.365 95.455 74.535 ;
        RECT 95.745 74.365 95.915 74.535 ;
        RECT 96.205 74.365 96.375 74.535 ;
        RECT 96.665 74.365 96.835 74.535 ;
        RECT 97.125 74.365 97.295 74.535 ;
        RECT 97.585 74.365 97.755 74.535 ;
        RECT 98.045 74.365 98.215 74.535 ;
        RECT 98.505 74.365 98.675 74.535 ;
        RECT 98.965 74.365 99.135 74.535 ;
        RECT 99.425 74.365 99.595 74.535 ;
        RECT 99.885 74.365 100.055 74.535 ;
        RECT 100.345 74.365 100.515 74.535 ;
        RECT 100.805 74.365 100.975 74.535 ;
        RECT 101.265 74.365 101.435 74.535 ;
        RECT 101.725 74.365 101.895 74.535 ;
        RECT 102.185 74.365 102.355 74.535 ;
        RECT 102.645 74.365 102.815 74.535 ;
        RECT 103.105 74.365 103.275 74.535 ;
        RECT 103.565 74.365 103.735 74.535 ;
        RECT 104.025 74.365 104.195 74.535 ;
        RECT 104.485 74.365 104.655 74.535 ;
        RECT 104.945 74.365 105.115 74.535 ;
        RECT 105.405 74.365 105.575 74.535 ;
        RECT 105.865 74.365 106.035 74.535 ;
        RECT 106.325 74.365 106.495 74.535 ;
        RECT 106.785 74.365 106.955 74.535 ;
        RECT 107.245 74.365 107.415 74.535 ;
        RECT 107.705 74.365 107.875 74.535 ;
        RECT 108.165 74.365 108.335 74.535 ;
        RECT 108.625 74.365 108.795 74.535 ;
        RECT 109.085 74.365 109.255 74.535 ;
        RECT 109.545 74.365 109.715 74.535 ;
        RECT 110.005 74.365 110.175 74.535 ;
        RECT 110.465 74.365 110.635 74.535 ;
        RECT 110.925 74.365 111.095 74.535 ;
        RECT 111.385 74.365 111.555 74.535 ;
        RECT 111.845 74.365 112.015 74.535 ;
        RECT 112.305 74.365 112.475 74.535 ;
        RECT 112.765 74.365 112.935 74.535 ;
        RECT 113.225 74.365 113.395 74.535 ;
        RECT 113.685 74.365 113.855 74.535 ;
        RECT 114.145 74.365 114.315 74.535 ;
        RECT 114.605 74.365 114.775 74.535 ;
        RECT 115.065 74.365 115.235 74.535 ;
        RECT 115.525 74.365 115.695 74.535 ;
        RECT 115.985 74.365 116.155 74.535 ;
        RECT 116.445 74.365 116.615 74.535 ;
        RECT 116.905 74.365 117.075 74.535 ;
        RECT 117.365 74.365 117.535 74.535 ;
        RECT 117.825 74.365 117.995 74.535 ;
        RECT 118.285 74.365 118.455 74.535 ;
        RECT 118.745 74.365 118.915 74.535 ;
        RECT 119.205 74.365 119.375 74.535 ;
        RECT 119.665 74.365 119.835 74.535 ;
        RECT 120.125 74.365 120.295 74.535 ;
        RECT 120.585 74.365 120.755 74.535 ;
        RECT 121.045 74.365 121.215 74.535 ;
        RECT 121.505 74.365 121.675 74.535 ;
        RECT 121.965 74.365 122.135 74.535 ;
        RECT 122.425 74.365 122.595 74.535 ;
        RECT 122.885 74.365 123.055 74.535 ;
        RECT 123.345 74.365 123.515 74.535 ;
        RECT 123.805 74.365 123.975 74.535 ;
        RECT 124.265 74.365 124.435 74.535 ;
        RECT 124.725 74.365 124.895 74.535 ;
        RECT 125.185 74.365 125.355 74.535 ;
        RECT 125.645 74.365 125.815 74.535 ;
        RECT 126.105 74.365 126.275 74.535 ;
        RECT 126.565 74.365 126.735 74.535 ;
        RECT 127.025 74.365 127.195 74.535 ;
        RECT 127.485 74.365 127.655 74.535 ;
        RECT 127.945 74.365 128.115 74.535 ;
        RECT 128.405 74.365 128.575 74.535 ;
        RECT 128.865 74.365 129.035 74.535 ;
        RECT 129.325 74.365 129.495 74.535 ;
        RECT 129.785 74.365 129.955 74.535 ;
        RECT 130.245 74.365 130.415 74.535 ;
        RECT 130.705 74.365 130.875 74.535 ;
        RECT 131.165 74.365 131.335 74.535 ;
        RECT 131.625 74.365 131.795 74.535 ;
        RECT 132.085 74.365 132.255 74.535 ;
        RECT 132.545 74.365 132.715 74.535 ;
        RECT 133.005 74.365 133.175 74.535 ;
        RECT 133.465 74.365 133.635 74.535 ;
        RECT 133.925 74.365 134.095 74.535 ;
        RECT 134.385 74.365 134.555 74.535 ;
        RECT 134.845 74.365 135.015 74.535 ;
        RECT 135.305 74.365 135.475 74.535 ;
        RECT 135.765 74.365 135.935 74.535 ;
        RECT 136.225 74.365 136.395 74.535 ;
        RECT 136.685 74.365 136.855 74.535 ;
        RECT 137.145 74.365 137.315 74.535 ;
        RECT 137.605 74.365 137.775 74.535 ;
        RECT 138.065 74.365 138.235 74.535 ;
        RECT 138.525 74.365 138.695 74.535 ;
        RECT 138.985 74.365 139.155 74.535 ;
        RECT 50.665 71.645 50.835 71.815 ;
        RECT 51.125 71.645 51.295 71.815 ;
        RECT 51.585 71.645 51.755 71.815 ;
        RECT 52.045 71.645 52.215 71.815 ;
        RECT 52.505 71.645 52.675 71.815 ;
        RECT 52.965 71.645 53.135 71.815 ;
        RECT 53.425 71.645 53.595 71.815 ;
        RECT 53.885 71.645 54.055 71.815 ;
        RECT 54.345 71.645 54.515 71.815 ;
        RECT 54.805 71.645 54.975 71.815 ;
        RECT 55.265 71.645 55.435 71.815 ;
        RECT 55.725 71.645 55.895 71.815 ;
        RECT 56.185 71.645 56.355 71.815 ;
        RECT 56.645 71.645 56.815 71.815 ;
        RECT 57.105 71.645 57.275 71.815 ;
        RECT 57.565 71.645 57.735 71.815 ;
        RECT 58.025 71.645 58.195 71.815 ;
        RECT 58.485 71.645 58.655 71.815 ;
        RECT 58.945 71.645 59.115 71.815 ;
        RECT 59.405 71.645 59.575 71.815 ;
        RECT 59.865 71.645 60.035 71.815 ;
        RECT 60.325 71.645 60.495 71.815 ;
        RECT 60.785 71.645 60.955 71.815 ;
        RECT 61.245 71.645 61.415 71.815 ;
        RECT 61.705 71.645 61.875 71.815 ;
        RECT 62.165 71.645 62.335 71.815 ;
        RECT 62.625 71.645 62.795 71.815 ;
        RECT 63.085 71.645 63.255 71.815 ;
        RECT 63.545 71.645 63.715 71.815 ;
        RECT 64.005 71.645 64.175 71.815 ;
        RECT 64.465 71.645 64.635 71.815 ;
        RECT 64.925 71.645 65.095 71.815 ;
        RECT 65.385 71.645 65.555 71.815 ;
        RECT 65.845 71.645 66.015 71.815 ;
        RECT 66.305 71.645 66.475 71.815 ;
        RECT 66.765 71.645 66.935 71.815 ;
        RECT 67.225 71.645 67.395 71.815 ;
        RECT 67.685 71.645 67.855 71.815 ;
        RECT 68.145 71.645 68.315 71.815 ;
        RECT 68.605 71.645 68.775 71.815 ;
        RECT 69.065 71.645 69.235 71.815 ;
        RECT 69.525 71.645 69.695 71.815 ;
        RECT 69.985 71.645 70.155 71.815 ;
        RECT 70.445 71.645 70.615 71.815 ;
        RECT 70.905 71.645 71.075 71.815 ;
        RECT 71.365 71.645 71.535 71.815 ;
        RECT 71.825 71.645 71.995 71.815 ;
        RECT 72.285 71.645 72.455 71.815 ;
        RECT 72.745 71.645 72.915 71.815 ;
        RECT 73.205 71.645 73.375 71.815 ;
        RECT 73.665 71.645 73.835 71.815 ;
        RECT 74.125 71.645 74.295 71.815 ;
        RECT 74.585 71.645 74.755 71.815 ;
        RECT 75.045 71.645 75.215 71.815 ;
        RECT 75.505 71.645 75.675 71.815 ;
        RECT 75.965 71.645 76.135 71.815 ;
        RECT 76.425 71.645 76.595 71.815 ;
        RECT 76.885 71.645 77.055 71.815 ;
        RECT 77.345 71.645 77.515 71.815 ;
        RECT 77.805 71.645 77.975 71.815 ;
        RECT 78.265 71.645 78.435 71.815 ;
        RECT 78.725 71.645 78.895 71.815 ;
        RECT 79.185 71.645 79.355 71.815 ;
        RECT 79.645 71.645 79.815 71.815 ;
        RECT 80.105 71.645 80.275 71.815 ;
        RECT 80.565 71.645 80.735 71.815 ;
        RECT 81.025 71.645 81.195 71.815 ;
        RECT 81.485 71.645 81.655 71.815 ;
        RECT 81.945 71.645 82.115 71.815 ;
        RECT 82.405 71.645 82.575 71.815 ;
        RECT 82.865 71.645 83.035 71.815 ;
        RECT 83.325 71.645 83.495 71.815 ;
        RECT 83.785 71.645 83.955 71.815 ;
        RECT 84.245 71.645 84.415 71.815 ;
        RECT 84.705 71.645 84.875 71.815 ;
        RECT 85.165 71.645 85.335 71.815 ;
        RECT 85.625 71.645 85.795 71.815 ;
        RECT 86.085 71.645 86.255 71.815 ;
        RECT 86.545 71.645 86.715 71.815 ;
        RECT 87.005 71.645 87.175 71.815 ;
        RECT 87.465 71.645 87.635 71.815 ;
        RECT 87.925 71.645 88.095 71.815 ;
        RECT 88.385 71.645 88.555 71.815 ;
        RECT 88.845 71.645 89.015 71.815 ;
        RECT 89.305 71.645 89.475 71.815 ;
        RECT 89.765 71.645 89.935 71.815 ;
        RECT 90.225 71.645 90.395 71.815 ;
        RECT 90.685 71.645 90.855 71.815 ;
        RECT 91.145 71.645 91.315 71.815 ;
        RECT 91.605 71.645 91.775 71.815 ;
        RECT 92.065 71.645 92.235 71.815 ;
        RECT 92.525 71.645 92.695 71.815 ;
        RECT 92.985 71.645 93.155 71.815 ;
        RECT 93.445 71.645 93.615 71.815 ;
        RECT 93.905 71.645 94.075 71.815 ;
        RECT 94.365 71.645 94.535 71.815 ;
        RECT 94.825 71.645 94.995 71.815 ;
        RECT 95.285 71.645 95.455 71.815 ;
        RECT 95.745 71.645 95.915 71.815 ;
        RECT 96.205 71.645 96.375 71.815 ;
        RECT 96.665 71.645 96.835 71.815 ;
        RECT 97.125 71.645 97.295 71.815 ;
        RECT 97.585 71.645 97.755 71.815 ;
        RECT 98.045 71.645 98.215 71.815 ;
        RECT 98.505 71.645 98.675 71.815 ;
        RECT 98.965 71.645 99.135 71.815 ;
        RECT 99.425 71.645 99.595 71.815 ;
        RECT 99.885 71.645 100.055 71.815 ;
        RECT 100.345 71.645 100.515 71.815 ;
        RECT 100.805 71.645 100.975 71.815 ;
        RECT 101.265 71.645 101.435 71.815 ;
        RECT 101.725 71.645 101.895 71.815 ;
        RECT 102.185 71.645 102.355 71.815 ;
        RECT 102.645 71.645 102.815 71.815 ;
        RECT 103.105 71.645 103.275 71.815 ;
        RECT 103.565 71.645 103.735 71.815 ;
        RECT 104.025 71.645 104.195 71.815 ;
        RECT 104.485 71.645 104.655 71.815 ;
        RECT 104.945 71.645 105.115 71.815 ;
        RECT 105.405 71.645 105.575 71.815 ;
        RECT 105.865 71.645 106.035 71.815 ;
        RECT 106.325 71.645 106.495 71.815 ;
        RECT 106.785 71.645 106.955 71.815 ;
        RECT 107.245 71.645 107.415 71.815 ;
        RECT 107.705 71.645 107.875 71.815 ;
        RECT 108.165 71.645 108.335 71.815 ;
        RECT 108.625 71.645 108.795 71.815 ;
        RECT 109.085 71.645 109.255 71.815 ;
        RECT 109.545 71.645 109.715 71.815 ;
        RECT 110.005 71.645 110.175 71.815 ;
        RECT 110.465 71.645 110.635 71.815 ;
        RECT 110.925 71.645 111.095 71.815 ;
        RECT 111.385 71.645 111.555 71.815 ;
        RECT 111.845 71.645 112.015 71.815 ;
        RECT 112.305 71.645 112.475 71.815 ;
        RECT 112.765 71.645 112.935 71.815 ;
        RECT 113.225 71.645 113.395 71.815 ;
        RECT 113.685 71.645 113.855 71.815 ;
        RECT 114.145 71.645 114.315 71.815 ;
        RECT 114.605 71.645 114.775 71.815 ;
        RECT 115.065 71.645 115.235 71.815 ;
        RECT 115.525 71.645 115.695 71.815 ;
        RECT 115.985 71.645 116.155 71.815 ;
        RECT 116.445 71.645 116.615 71.815 ;
        RECT 116.905 71.645 117.075 71.815 ;
        RECT 117.365 71.645 117.535 71.815 ;
        RECT 117.825 71.645 117.995 71.815 ;
        RECT 118.285 71.645 118.455 71.815 ;
        RECT 118.745 71.645 118.915 71.815 ;
        RECT 119.205 71.645 119.375 71.815 ;
        RECT 119.665 71.645 119.835 71.815 ;
        RECT 120.125 71.645 120.295 71.815 ;
        RECT 120.585 71.645 120.755 71.815 ;
        RECT 121.045 71.645 121.215 71.815 ;
        RECT 121.505 71.645 121.675 71.815 ;
        RECT 121.965 71.645 122.135 71.815 ;
        RECT 122.425 71.645 122.595 71.815 ;
        RECT 122.885 71.645 123.055 71.815 ;
        RECT 123.345 71.645 123.515 71.815 ;
        RECT 123.805 71.645 123.975 71.815 ;
        RECT 124.265 71.645 124.435 71.815 ;
        RECT 124.725 71.645 124.895 71.815 ;
        RECT 125.185 71.645 125.355 71.815 ;
        RECT 125.645 71.645 125.815 71.815 ;
        RECT 126.105 71.645 126.275 71.815 ;
        RECT 126.565 71.645 126.735 71.815 ;
        RECT 127.025 71.645 127.195 71.815 ;
        RECT 127.485 71.645 127.655 71.815 ;
        RECT 127.945 71.645 128.115 71.815 ;
        RECT 128.405 71.645 128.575 71.815 ;
        RECT 128.865 71.645 129.035 71.815 ;
        RECT 129.325 71.645 129.495 71.815 ;
        RECT 129.785 71.645 129.955 71.815 ;
        RECT 130.245 71.645 130.415 71.815 ;
        RECT 130.705 71.645 130.875 71.815 ;
        RECT 131.165 71.645 131.335 71.815 ;
        RECT 131.625 71.645 131.795 71.815 ;
        RECT 132.085 71.645 132.255 71.815 ;
        RECT 132.545 71.645 132.715 71.815 ;
        RECT 133.005 71.645 133.175 71.815 ;
        RECT 133.465 71.645 133.635 71.815 ;
        RECT 133.925 71.645 134.095 71.815 ;
        RECT 134.385 71.645 134.555 71.815 ;
        RECT 134.845 71.645 135.015 71.815 ;
        RECT 135.305 71.645 135.475 71.815 ;
        RECT 135.765 71.645 135.935 71.815 ;
        RECT 136.225 71.645 136.395 71.815 ;
        RECT 136.685 71.645 136.855 71.815 ;
        RECT 137.145 71.645 137.315 71.815 ;
        RECT 137.605 71.645 137.775 71.815 ;
        RECT 138.065 71.645 138.235 71.815 ;
        RECT 138.525 71.645 138.695 71.815 ;
        RECT 138.985 71.645 139.155 71.815 ;
        RECT 50.665 68.925 50.835 69.095 ;
        RECT 51.125 68.925 51.295 69.095 ;
        RECT 51.585 68.925 51.755 69.095 ;
        RECT 52.045 68.925 52.215 69.095 ;
        RECT 52.505 68.925 52.675 69.095 ;
        RECT 52.965 68.925 53.135 69.095 ;
        RECT 53.425 68.925 53.595 69.095 ;
        RECT 53.885 68.925 54.055 69.095 ;
        RECT 54.345 68.925 54.515 69.095 ;
        RECT 54.805 68.925 54.975 69.095 ;
        RECT 55.265 68.925 55.435 69.095 ;
        RECT 55.725 68.925 55.895 69.095 ;
        RECT 56.185 68.925 56.355 69.095 ;
        RECT 56.645 68.925 56.815 69.095 ;
        RECT 57.105 68.925 57.275 69.095 ;
        RECT 57.565 68.925 57.735 69.095 ;
        RECT 58.025 68.925 58.195 69.095 ;
        RECT 58.485 68.925 58.655 69.095 ;
        RECT 58.945 68.925 59.115 69.095 ;
        RECT 59.405 68.925 59.575 69.095 ;
        RECT 59.865 68.925 60.035 69.095 ;
        RECT 60.325 68.925 60.495 69.095 ;
        RECT 60.785 68.925 60.955 69.095 ;
        RECT 61.245 68.925 61.415 69.095 ;
        RECT 61.705 68.925 61.875 69.095 ;
        RECT 62.165 68.925 62.335 69.095 ;
        RECT 62.625 68.925 62.795 69.095 ;
        RECT 63.085 68.925 63.255 69.095 ;
        RECT 63.545 68.925 63.715 69.095 ;
        RECT 64.005 68.925 64.175 69.095 ;
        RECT 64.465 68.925 64.635 69.095 ;
        RECT 64.925 68.925 65.095 69.095 ;
        RECT 65.385 68.925 65.555 69.095 ;
        RECT 65.845 68.925 66.015 69.095 ;
        RECT 66.305 68.925 66.475 69.095 ;
        RECT 66.765 68.925 66.935 69.095 ;
        RECT 67.225 68.925 67.395 69.095 ;
        RECT 67.685 68.925 67.855 69.095 ;
        RECT 68.145 68.925 68.315 69.095 ;
        RECT 68.605 68.925 68.775 69.095 ;
        RECT 69.065 68.925 69.235 69.095 ;
        RECT 69.525 68.925 69.695 69.095 ;
        RECT 69.985 68.925 70.155 69.095 ;
        RECT 70.445 68.925 70.615 69.095 ;
        RECT 70.905 68.925 71.075 69.095 ;
        RECT 71.365 68.925 71.535 69.095 ;
        RECT 71.825 68.925 71.995 69.095 ;
        RECT 72.285 68.925 72.455 69.095 ;
        RECT 72.745 68.925 72.915 69.095 ;
        RECT 73.205 68.925 73.375 69.095 ;
        RECT 73.665 68.925 73.835 69.095 ;
        RECT 74.125 68.925 74.295 69.095 ;
        RECT 74.585 68.925 74.755 69.095 ;
        RECT 75.045 68.925 75.215 69.095 ;
        RECT 75.505 68.925 75.675 69.095 ;
        RECT 75.965 68.925 76.135 69.095 ;
        RECT 76.425 68.925 76.595 69.095 ;
        RECT 76.885 68.925 77.055 69.095 ;
        RECT 77.345 68.925 77.515 69.095 ;
        RECT 77.805 68.925 77.975 69.095 ;
        RECT 78.265 68.925 78.435 69.095 ;
        RECT 78.725 68.925 78.895 69.095 ;
        RECT 79.185 68.925 79.355 69.095 ;
        RECT 79.645 68.925 79.815 69.095 ;
        RECT 80.105 68.925 80.275 69.095 ;
        RECT 80.565 68.925 80.735 69.095 ;
        RECT 81.025 68.925 81.195 69.095 ;
        RECT 81.485 68.925 81.655 69.095 ;
        RECT 81.945 68.925 82.115 69.095 ;
        RECT 82.405 68.925 82.575 69.095 ;
        RECT 82.865 68.925 83.035 69.095 ;
        RECT 83.325 68.925 83.495 69.095 ;
        RECT 83.785 68.925 83.955 69.095 ;
        RECT 84.245 68.925 84.415 69.095 ;
        RECT 84.705 68.925 84.875 69.095 ;
        RECT 85.165 68.925 85.335 69.095 ;
        RECT 85.625 68.925 85.795 69.095 ;
        RECT 86.085 68.925 86.255 69.095 ;
        RECT 86.545 68.925 86.715 69.095 ;
        RECT 87.005 68.925 87.175 69.095 ;
        RECT 87.465 68.925 87.635 69.095 ;
        RECT 87.925 68.925 88.095 69.095 ;
        RECT 88.385 68.925 88.555 69.095 ;
        RECT 88.845 68.925 89.015 69.095 ;
        RECT 89.305 68.925 89.475 69.095 ;
        RECT 89.765 68.925 89.935 69.095 ;
        RECT 90.225 68.925 90.395 69.095 ;
        RECT 90.685 68.925 90.855 69.095 ;
        RECT 91.145 68.925 91.315 69.095 ;
        RECT 91.605 68.925 91.775 69.095 ;
        RECT 92.065 68.925 92.235 69.095 ;
        RECT 92.525 68.925 92.695 69.095 ;
        RECT 92.985 68.925 93.155 69.095 ;
        RECT 93.445 68.925 93.615 69.095 ;
        RECT 93.905 68.925 94.075 69.095 ;
        RECT 94.365 68.925 94.535 69.095 ;
        RECT 94.825 68.925 94.995 69.095 ;
        RECT 95.285 68.925 95.455 69.095 ;
        RECT 95.745 68.925 95.915 69.095 ;
        RECT 96.205 68.925 96.375 69.095 ;
        RECT 96.665 68.925 96.835 69.095 ;
        RECT 97.125 68.925 97.295 69.095 ;
        RECT 97.585 68.925 97.755 69.095 ;
        RECT 98.045 68.925 98.215 69.095 ;
        RECT 98.505 68.925 98.675 69.095 ;
        RECT 98.965 68.925 99.135 69.095 ;
        RECT 99.425 68.925 99.595 69.095 ;
        RECT 99.885 68.925 100.055 69.095 ;
        RECT 100.345 68.925 100.515 69.095 ;
        RECT 100.805 68.925 100.975 69.095 ;
        RECT 101.265 68.925 101.435 69.095 ;
        RECT 101.725 68.925 101.895 69.095 ;
        RECT 102.185 68.925 102.355 69.095 ;
        RECT 102.645 68.925 102.815 69.095 ;
        RECT 103.105 68.925 103.275 69.095 ;
        RECT 103.565 68.925 103.735 69.095 ;
        RECT 104.025 68.925 104.195 69.095 ;
        RECT 104.485 68.925 104.655 69.095 ;
        RECT 104.945 68.925 105.115 69.095 ;
        RECT 105.405 68.925 105.575 69.095 ;
        RECT 105.865 68.925 106.035 69.095 ;
        RECT 106.325 68.925 106.495 69.095 ;
        RECT 106.785 68.925 106.955 69.095 ;
        RECT 107.245 68.925 107.415 69.095 ;
        RECT 107.705 68.925 107.875 69.095 ;
        RECT 108.165 68.925 108.335 69.095 ;
        RECT 108.625 68.925 108.795 69.095 ;
        RECT 109.085 68.925 109.255 69.095 ;
        RECT 109.545 68.925 109.715 69.095 ;
        RECT 110.005 68.925 110.175 69.095 ;
        RECT 110.465 68.925 110.635 69.095 ;
        RECT 110.925 68.925 111.095 69.095 ;
        RECT 111.385 68.925 111.555 69.095 ;
        RECT 111.845 68.925 112.015 69.095 ;
        RECT 112.305 68.925 112.475 69.095 ;
        RECT 112.765 68.925 112.935 69.095 ;
        RECT 113.225 68.925 113.395 69.095 ;
        RECT 113.685 68.925 113.855 69.095 ;
        RECT 114.145 68.925 114.315 69.095 ;
        RECT 114.605 68.925 114.775 69.095 ;
        RECT 115.065 68.925 115.235 69.095 ;
        RECT 115.525 68.925 115.695 69.095 ;
        RECT 115.985 68.925 116.155 69.095 ;
        RECT 116.445 68.925 116.615 69.095 ;
        RECT 116.905 68.925 117.075 69.095 ;
        RECT 117.365 68.925 117.535 69.095 ;
        RECT 117.825 68.925 117.995 69.095 ;
        RECT 118.285 68.925 118.455 69.095 ;
        RECT 118.745 68.925 118.915 69.095 ;
        RECT 119.205 68.925 119.375 69.095 ;
        RECT 119.665 68.925 119.835 69.095 ;
        RECT 120.125 68.925 120.295 69.095 ;
        RECT 120.585 68.925 120.755 69.095 ;
        RECT 121.045 68.925 121.215 69.095 ;
        RECT 121.505 68.925 121.675 69.095 ;
        RECT 121.965 68.925 122.135 69.095 ;
        RECT 122.425 68.925 122.595 69.095 ;
        RECT 122.885 68.925 123.055 69.095 ;
        RECT 123.345 68.925 123.515 69.095 ;
        RECT 123.805 68.925 123.975 69.095 ;
        RECT 124.265 68.925 124.435 69.095 ;
        RECT 124.725 68.925 124.895 69.095 ;
        RECT 125.185 68.925 125.355 69.095 ;
        RECT 125.645 68.925 125.815 69.095 ;
        RECT 126.105 68.925 126.275 69.095 ;
        RECT 126.565 68.925 126.735 69.095 ;
        RECT 127.025 68.925 127.195 69.095 ;
        RECT 127.485 68.925 127.655 69.095 ;
        RECT 127.945 68.925 128.115 69.095 ;
        RECT 128.405 68.925 128.575 69.095 ;
        RECT 128.865 68.925 129.035 69.095 ;
        RECT 129.325 68.925 129.495 69.095 ;
        RECT 129.785 68.925 129.955 69.095 ;
        RECT 130.245 68.925 130.415 69.095 ;
        RECT 130.705 68.925 130.875 69.095 ;
        RECT 131.165 68.925 131.335 69.095 ;
        RECT 131.625 68.925 131.795 69.095 ;
        RECT 132.085 68.925 132.255 69.095 ;
        RECT 132.545 68.925 132.715 69.095 ;
        RECT 133.005 68.925 133.175 69.095 ;
        RECT 133.465 68.925 133.635 69.095 ;
        RECT 133.925 68.925 134.095 69.095 ;
        RECT 134.385 68.925 134.555 69.095 ;
        RECT 134.845 68.925 135.015 69.095 ;
        RECT 135.305 68.925 135.475 69.095 ;
        RECT 135.765 68.925 135.935 69.095 ;
        RECT 136.225 68.925 136.395 69.095 ;
        RECT 136.685 68.925 136.855 69.095 ;
        RECT 137.145 68.925 137.315 69.095 ;
        RECT 137.605 68.925 137.775 69.095 ;
        RECT 138.065 68.925 138.235 69.095 ;
        RECT 138.525 68.925 138.695 69.095 ;
        RECT 138.985 68.925 139.155 69.095 ;
        RECT 50.665 66.205 50.835 66.375 ;
        RECT 51.125 66.205 51.295 66.375 ;
        RECT 51.585 66.205 51.755 66.375 ;
        RECT 52.045 66.205 52.215 66.375 ;
        RECT 52.505 66.205 52.675 66.375 ;
        RECT 52.965 66.205 53.135 66.375 ;
        RECT 53.425 66.205 53.595 66.375 ;
        RECT 53.885 66.205 54.055 66.375 ;
        RECT 54.345 66.205 54.515 66.375 ;
        RECT 54.805 66.205 54.975 66.375 ;
        RECT 55.265 66.205 55.435 66.375 ;
        RECT 55.725 66.205 55.895 66.375 ;
        RECT 56.185 66.205 56.355 66.375 ;
        RECT 56.645 66.205 56.815 66.375 ;
        RECT 57.105 66.205 57.275 66.375 ;
        RECT 57.565 66.205 57.735 66.375 ;
        RECT 58.025 66.205 58.195 66.375 ;
        RECT 58.485 66.205 58.655 66.375 ;
        RECT 58.945 66.205 59.115 66.375 ;
        RECT 59.405 66.205 59.575 66.375 ;
        RECT 59.865 66.205 60.035 66.375 ;
        RECT 60.325 66.205 60.495 66.375 ;
        RECT 60.785 66.205 60.955 66.375 ;
        RECT 61.245 66.205 61.415 66.375 ;
        RECT 61.705 66.205 61.875 66.375 ;
        RECT 62.165 66.205 62.335 66.375 ;
        RECT 62.625 66.205 62.795 66.375 ;
        RECT 63.085 66.205 63.255 66.375 ;
        RECT 63.545 66.205 63.715 66.375 ;
        RECT 64.005 66.205 64.175 66.375 ;
        RECT 64.465 66.205 64.635 66.375 ;
        RECT 64.925 66.205 65.095 66.375 ;
        RECT 65.385 66.205 65.555 66.375 ;
        RECT 65.845 66.205 66.015 66.375 ;
        RECT 66.305 66.205 66.475 66.375 ;
        RECT 66.765 66.205 66.935 66.375 ;
        RECT 67.225 66.205 67.395 66.375 ;
        RECT 67.685 66.205 67.855 66.375 ;
        RECT 68.145 66.205 68.315 66.375 ;
        RECT 68.605 66.205 68.775 66.375 ;
        RECT 69.065 66.205 69.235 66.375 ;
        RECT 69.525 66.205 69.695 66.375 ;
        RECT 69.985 66.205 70.155 66.375 ;
        RECT 70.445 66.205 70.615 66.375 ;
        RECT 70.905 66.205 71.075 66.375 ;
        RECT 71.365 66.205 71.535 66.375 ;
        RECT 71.825 66.205 71.995 66.375 ;
        RECT 72.285 66.205 72.455 66.375 ;
        RECT 72.745 66.205 72.915 66.375 ;
        RECT 73.205 66.205 73.375 66.375 ;
        RECT 73.665 66.205 73.835 66.375 ;
        RECT 74.125 66.205 74.295 66.375 ;
        RECT 74.585 66.205 74.755 66.375 ;
        RECT 75.045 66.205 75.215 66.375 ;
        RECT 75.505 66.205 75.675 66.375 ;
        RECT 75.965 66.205 76.135 66.375 ;
        RECT 76.425 66.205 76.595 66.375 ;
        RECT 76.885 66.205 77.055 66.375 ;
        RECT 77.345 66.205 77.515 66.375 ;
        RECT 77.805 66.205 77.975 66.375 ;
        RECT 78.265 66.205 78.435 66.375 ;
        RECT 78.725 66.205 78.895 66.375 ;
        RECT 79.185 66.205 79.355 66.375 ;
        RECT 79.645 66.205 79.815 66.375 ;
        RECT 80.105 66.205 80.275 66.375 ;
        RECT 80.565 66.205 80.735 66.375 ;
        RECT 81.025 66.205 81.195 66.375 ;
        RECT 81.485 66.205 81.655 66.375 ;
        RECT 81.945 66.205 82.115 66.375 ;
        RECT 82.405 66.205 82.575 66.375 ;
        RECT 82.865 66.205 83.035 66.375 ;
        RECT 83.325 66.205 83.495 66.375 ;
        RECT 83.785 66.205 83.955 66.375 ;
        RECT 84.245 66.205 84.415 66.375 ;
        RECT 84.705 66.205 84.875 66.375 ;
        RECT 85.165 66.205 85.335 66.375 ;
        RECT 85.625 66.205 85.795 66.375 ;
        RECT 86.085 66.205 86.255 66.375 ;
        RECT 86.545 66.205 86.715 66.375 ;
        RECT 87.005 66.205 87.175 66.375 ;
        RECT 87.465 66.205 87.635 66.375 ;
        RECT 87.925 66.205 88.095 66.375 ;
        RECT 88.385 66.205 88.555 66.375 ;
        RECT 88.845 66.205 89.015 66.375 ;
        RECT 89.305 66.205 89.475 66.375 ;
        RECT 89.765 66.205 89.935 66.375 ;
        RECT 90.225 66.205 90.395 66.375 ;
        RECT 90.685 66.205 90.855 66.375 ;
        RECT 91.145 66.205 91.315 66.375 ;
        RECT 91.605 66.205 91.775 66.375 ;
        RECT 92.065 66.205 92.235 66.375 ;
        RECT 92.525 66.205 92.695 66.375 ;
        RECT 92.985 66.205 93.155 66.375 ;
        RECT 93.445 66.205 93.615 66.375 ;
        RECT 93.905 66.205 94.075 66.375 ;
        RECT 94.365 66.205 94.535 66.375 ;
        RECT 94.825 66.205 94.995 66.375 ;
        RECT 95.285 66.205 95.455 66.375 ;
        RECT 95.745 66.205 95.915 66.375 ;
        RECT 96.205 66.205 96.375 66.375 ;
        RECT 96.665 66.205 96.835 66.375 ;
        RECT 97.125 66.205 97.295 66.375 ;
        RECT 97.585 66.205 97.755 66.375 ;
        RECT 98.045 66.205 98.215 66.375 ;
        RECT 98.505 66.205 98.675 66.375 ;
        RECT 98.965 66.205 99.135 66.375 ;
        RECT 99.425 66.205 99.595 66.375 ;
        RECT 99.885 66.205 100.055 66.375 ;
        RECT 100.345 66.205 100.515 66.375 ;
        RECT 100.805 66.205 100.975 66.375 ;
        RECT 101.265 66.205 101.435 66.375 ;
        RECT 101.725 66.205 101.895 66.375 ;
        RECT 102.185 66.205 102.355 66.375 ;
        RECT 102.645 66.205 102.815 66.375 ;
        RECT 103.105 66.205 103.275 66.375 ;
        RECT 103.565 66.205 103.735 66.375 ;
        RECT 104.025 66.205 104.195 66.375 ;
        RECT 104.485 66.205 104.655 66.375 ;
        RECT 104.945 66.205 105.115 66.375 ;
        RECT 105.405 66.205 105.575 66.375 ;
        RECT 105.865 66.205 106.035 66.375 ;
        RECT 106.325 66.205 106.495 66.375 ;
        RECT 106.785 66.205 106.955 66.375 ;
        RECT 107.245 66.205 107.415 66.375 ;
        RECT 107.705 66.205 107.875 66.375 ;
        RECT 108.165 66.205 108.335 66.375 ;
        RECT 108.625 66.205 108.795 66.375 ;
        RECT 109.085 66.205 109.255 66.375 ;
        RECT 109.545 66.205 109.715 66.375 ;
        RECT 110.005 66.205 110.175 66.375 ;
        RECT 110.465 66.205 110.635 66.375 ;
        RECT 110.925 66.205 111.095 66.375 ;
        RECT 111.385 66.205 111.555 66.375 ;
        RECT 111.845 66.205 112.015 66.375 ;
        RECT 112.305 66.205 112.475 66.375 ;
        RECT 112.765 66.205 112.935 66.375 ;
        RECT 113.225 66.205 113.395 66.375 ;
        RECT 113.685 66.205 113.855 66.375 ;
        RECT 114.145 66.205 114.315 66.375 ;
        RECT 114.605 66.205 114.775 66.375 ;
        RECT 115.065 66.205 115.235 66.375 ;
        RECT 115.525 66.205 115.695 66.375 ;
        RECT 115.985 66.205 116.155 66.375 ;
        RECT 116.445 66.205 116.615 66.375 ;
        RECT 116.905 66.205 117.075 66.375 ;
        RECT 117.365 66.205 117.535 66.375 ;
        RECT 117.825 66.205 117.995 66.375 ;
        RECT 118.285 66.205 118.455 66.375 ;
        RECT 118.745 66.205 118.915 66.375 ;
        RECT 119.205 66.205 119.375 66.375 ;
        RECT 119.665 66.205 119.835 66.375 ;
        RECT 120.125 66.205 120.295 66.375 ;
        RECT 120.585 66.205 120.755 66.375 ;
        RECT 121.045 66.205 121.215 66.375 ;
        RECT 121.505 66.205 121.675 66.375 ;
        RECT 121.965 66.205 122.135 66.375 ;
        RECT 122.425 66.205 122.595 66.375 ;
        RECT 122.885 66.205 123.055 66.375 ;
        RECT 123.345 66.205 123.515 66.375 ;
        RECT 123.805 66.205 123.975 66.375 ;
        RECT 124.265 66.205 124.435 66.375 ;
        RECT 124.725 66.205 124.895 66.375 ;
        RECT 125.185 66.205 125.355 66.375 ;
        RECT 125.645 66.205 125.815 66.375 ;
        RECT 126.105 66.205 126.275 66.375 ;
        RECT 126.565 66.205 126.735 66.375 ;
        RECT 127.025 66.205 127.195 66.375 ;
        RECT 127.485 66.205 127.655 66.375 ;
        RECT 127.945 66.205 128.115 66.375 ;
        RECT 128.405 66.205 128.575 66.375 ;
        RECT 128.865 66.205 129.035 66.375 ;
        RECT 129.325 66.205 129.495 66.375 ;
        RECT 129.785 66.205 129.955 66.375 ;
        RECT 130.245 66.205 130.415 66.375 ;
        RECT 130.705 66.205 130.875 66.375 ;
        RECT 131.165 66.205 131.335 66.375 ;
        RECT 131.625 66.205 131.795 66.375 ;
        RECT 132.085 66.205 132.255 66.375 ;
        RECT 132.545 66.205 132.715 66.375 ;
        RECT 133.005 66.205 133.175 66.375 ;
        RECT 133.465 66.205 133.635 66.375 ;
        RECT 133.925 66.205 134.095 66.375 ;
        RECT 134.385 66.205 134.555 66.375 ;
        RECT 134.845 66.205 135.015 66.375 ;
        RECT 135.305 66.205 135.475 66.375 ;
        RECT 135.765 66.205 135.935 66.375 ;
        RECT 136.225 66.205 136.395 66.375 ;
        RECT 136.685 66.205 136.855 66.375 ;
        RECT 137.145 66.205 137.315 66.375 ;
        RECT 137.605 66.205 137.775 66.375 ;
        RECT 138.065 66.205 138.235 66.375 ;
        RECT 138.525 66.205 138.695 66.375 ;
        RECT 138.985 66.205 139.155 66.375 ;
        RECT 50.665 63.485 50.835 63.655 ;
        RECT 51.125 63.485 51.295 63.655 ;
        RECT 51.585 63.485 51.755 63.655 ;
        RECT 52.045 63.485 52.215 63.655 ;
        RECT 52.505 63.485 52.675 63.655 ;
        RECT 52.965 63.485 53.135 63.655 ;
        RECT 53.425 63.485 53.595 63.655 ;
        RECT 53.885 63.485 54.055 63.655 ;
        RECT 54.345 63.485 54.515 63.655 ;
        RECT 54.805 63.485 54.975 63.655 ;
        RECT 55.265 63.485 55.435 63.655 ;
        RECT 55.725 63.485 55.895 63.655 ;
        RECT 56.185 63.485 56.355 63.655 ;
        RECT 56.645 63.485 56.815 63.655 ;
        RECT 57.105 63.485 57.275 63.655 ;
        RECT 57.565 63.485 57.735 63.655 ;
        RECT 58.025 63.485 58.195 63.655 ;
        RECT 58.485 63.485 58.655 63.655 ;
        RECT 58.945 63.485 59.115 63.655 ;
        RECT 59.405 63.485 59.575 63.655 ;
        RECT 59.865 63.485 60.035 63.655 ;
        RECT 60.325 63.485 60.495 63.655 ;
        RECT 60.785 63.485 60.955 63.655 ;
        RECT 61.245 63.485 61.415 63.655 ;
        RECT 61.705 63.485 61.875 63.655 ;
        RECT 62.165 63.485 62.335 63.655 ;
        RECT 62.625 63.485 62.795 63.655 ;
        RECT 63.085 63.485 63.255 63.655 ;
        RECT 63.545 63.485 63.715 63.655 ;
        RECT 64.005 63.485 64.175 63.655 ;
        RECT 64.465 63.485 64.635 63.655 ;
        RECT 64.925 63.485 65.095 63.655 ;
        RECT 65.385 63.485 65.555 63.655 ;
        RECT 65.845 63.485 66.015 63.655 ;
        RECT 66.305 63.485 66.475 63.655 ;
        RECT 66.765 63.485 66.935 63.655 ;
        RECT 67.225 63.485 67.395 63.655 ;
        RECT 67.685 63.485 67.855 63.655 ;
        RECT 68.145 63.485 68.315 63.655 ;
        RECT 68.605 63.485 68.775 63.655 ;
        RECT 69.065 63.485 69.235 63.655 ;
        RECT 69.525 63.485 69.695 63.655 ;
        RECT 69.985 63.485 70.155 63.655 ;
        RECT 70.445 63.485 70.615 63.655 ;
        RECT 70.905 63.485 71.075 63.655 ;
        RECT 71.365 63.485 71.535 63.655 ;
        RECT 71.825 63.485 71.995 63.655 ;
        RECT 72.285 63.485 72.455 63.655 ;
        RECT 72.745 63.485 72.915 63.655 ;
        RECT 73.205 63.485 73.375 63.655 ;
        RECT 73.665 63.485 73.835 63.655 ;
        RECT 74.125 63.485 74.295 63.655 ;
        RECT 74.585 63.485 74.755 63.655 ;
        RECT 75.045 63.485 75.215 63.655 ;
        RECT 75.505 63.485 75.675 63.655 ;
        RECT 75.965 63.485 76.135 63.655 ;
        RECT 76.425 63.485 76.595 63.655 ;
        RECT 76.885 63.485 77.055 63.655 ;
        RECT 77.345 63.485 77.515 63.655 ;
        RECT 77.805 63.485 77.975 63.655 ;
        RECT 78.265 63.485 78.435 63.655 ;
        RECT 78.725 63.485 78.895 63.655 ;
        RECT 79.185 63.485 79.355 63.655 ;
        RECT 79.645 63.485 79.815 63.655 ;
        RECT 80.105 63.485 80.275 63.655 ;
        RECT 80.565 63.485 80.735 63.655 ;
        RECT 81.025 63.485 81.195 63.655 ;
        RECT 81.485 63.485 81.655 63.655 ;
        RECT 81.945 63.485 82.115 63.655 ;
        RECT 82.405 63.485 82.575 63.655 ;
        RECT 82.865 63.485 83.035 63.655 ;
        RECT 83.325 63.485 83.495 63.655 ;
        RECT 83.785 63.485 83.955 63.655 ;
        RECT 84.245 63.485 84.415 63.655 ;
        RECT 84.705 63.485 84.875 63.655 ;
        RECT 85.165 63.485 85.335 63.655 ;
        RECT 85.625 63.485 85.795 63.655 ;
        RECT 86.085 63.485 86.255 63.655 ;
        RECT 86.545 63.485 86.715 63.655 ;
        RECT 87.005 63.485 87.175 63.655 ;
        RECT 87.465 63.485 87.635 63.655 ;
        RECT 87.925 63.485 88.095 63.655 ;
        RECT 88.385 63.485 88.555 63.655 ;
        RECT 88.845 63.485 89.015 63.655 ;
        RECT 89.305 63.485 89.475 63.655 ;
        RECT 89.765 63.485 89.935 63.655 ;
        RECT 90.225 63.485 90.395 63.655 ;
        RECT 90.685 63.485 90.855 63.655 ;
        RECT 91.145 63.485 91.315 63.655 ;
        RECT 91.605 63.485 91.775 63.655 ;
        RECT 92.065 63.485 92.235 63.655 ;
        RECT 92.525 63.485 92.695 63.655 ;
        RECT 92.985 63.485 93.155 63.655 ;
        RECT 93.445 63.485 93.615 63.655 ;
        RECT 93.905 63.485 94.075 63.655 ;
        RECT 94.365 63.485 94.535 63.655 ;
        RECT 94.825 63.485 94.995 63.655 ;
        RECT 95.285 63.485 95.455 63.655 ;
        RECT 95.745 63.485 95.915 63.655 ;
        RECT 96.205 63.485 96.375 63.655 ;
        RECT 96.665 63.485 96.835 63.655 ;
        RECT 97.125 63.485 97.295 63.655 ;
        RECT 97.585 63.485 97.755 63.655 ;
        RECT 98.045 63.485 98.215 63.655 ;
        RECT 98.505 63.485 98.675 63.655 ;
        RECT 98.965 63.485 99.135 63.655 ;
        RECT 99.425 63.485 99.595 63.655 ;
        RECT 99.885 63.485 100.055 63.655 ;
        RECT 100.345 63.485 100.515 63.655 ;
        RECT 100.805 63.485 100.975 63.655 ;
        RECT 101.265 63.485 101.435 63.655 ;
        RECT 101.725 63.485 101.895 63.655 ;
        RECT 102.185 63.485 102.355 63.655 ;
        RECT 102.645 63.485 102.815 63.655 ;
        RECT 103.105 63.485 103.275 63.655 ;
        RECT 103.565 63.485 103.735 63.655 ;
        RECT 104.025 63.485 104.195 63.655 ;
        RECT 104.485 63.485 104.655 63.655 ;
        RECT 104.945 63.485 105.115 63.655 ;
        RECT 105.405 63.485 105.575 63.655 ;
        RECT 105.865 63.485 106.035 63.655 ;
        RECT 106.325 63.485 106.495 63.655 ;
        RECT 106.785 63.485 106.955 63.655 ;
        RECT 107.245 63.485 107.415 63.655 ;
        RECT 107.705 63.485 107.875 63.655 ;
        RECT 108.165 63.485 108.335 63.655 ;
        RECT 108.625 63.485 108.795 63.655 ;
        RECT 109.085 63.485 109.255 63.655 ;
        RECT 109.545 63.485 109.715 63.655 ;
        RECT 110.005 63.485 110.175 63.655 ;
        RECT 110.465 63.485 110.635 63.655 ;
        RECT 110.925 63.485 111.095 63.655 ;
        RECT 111.385 63.485 111.555 63.655 ;
        RECT 111.845 63.485 112.015 63.655 ;
        RECT 112.305 63.485 112.475 63.655 ;
        RECT 112.765 63.485 112.935 63.655 ;
        RECT 113.225 63.485 113.395 63.655 ;
        RECT 113.685 63.485 113.855 63.655 ;
        RECT 114.145 63.485 114.315 63.655 ;
        RECT 114.605 63.485 114.775 63.655 ;
        RECT 115.065 63.485 115.235 63.655 ;
        RECT 115.525 63.485 115.695 63.655 ;
        RECT 115.985 63.485 116.155 63.655 ;
        RECT 116.445 63.485 116.615 63.655 ;
        RECT 116.905 63.485 117.075 63.655 ;
        RECT 117.365 63.485 117.535 63.655 ;
        RECT 117.825 63.485 117.995 63.655 ;
        RECT 118.285 63.485 118.455 63.655 ;
        RECT 118.745 63.485 118.915 63.655 ;
        RECT 119.205 63.485 119.375 63.655 ;
        RECT 119.665 63.485 119.835 63.655 ;
        RECT 120.125 63.485 120.295 63.655 ;
        RECT 120.585 63.485 120.755 63.655 ;
        RECT 121.045 63.485 121.215 63.655 ;
        RECT 121.505 63.485 121.675 63.655 ;
        RECT 121.965 63.485 122.135 63.655 ;
        RECT 122.425 63.485 122.595 63.655 ;
        RECT 122.885 63.485 123.055 63.655 ;
        RECT 123.345 63.485 123.515 63.655 ;
        RECT 123.805 63.485 123.975 63.655 ;
        RECT 124.265 63.485 124.435 63.655 ;
        RECT 124.725 63.485 124.895 63.655 ;
        RECT 125.185 63.485 125.355 63.655 ;
        RECT 125.645 63.485 125.815 63.655 ;
        RECT 126.105 63.485 126.275 63.655 ;
        RECT 126.565 63.485 126.735 63.655 ;
        RECT 127.025 63.485 127.195 63.655 ;
        RECT 127.485 63.485 127.655 63.655 ;
        RECT 127.945 63.485 128.115 63.655 ;
        RECT 128.405 63.485 128.575 63.655 ;
        RECT 128.865 63.485 129.035 63.655 ;
        RECT 129.325 63.485 129.495 63.655 ;
        RECT 129.785 63.485 129.955 63.655 ;
        RECT 130.245 63.485 130.415 63.655 ;
        RECT 130.705 63.485 130.875 63.655 ;
        RECT 131.165 63.485 131.335 63.655 ;
        RECT 131.625 63.485 131.795 63.655 ;
        RECT 132.085 63.485 132.255 63.655 ;
        RECT 132.545 63.485 132.715 63.655 ;
        RECT 133.005 63.485 133.175 63.655 ;
        RECT 133.465 63.485 133.635 63.655 ;
        RECT 133.925 63.485 134.095 63.655 ;
        RECT 134.385 63.485 134.555 63.655 ;
        RECT 134.845 63.485 135.015 63.655 ;
        RECT 135.305 63.485 135.475 63.655 ;
        RECT 135.765 63.485 135.935 63.655 ;
        RECT 136.225 63.485 136.395 63.655 ;
        RECT 136.685 63.485 136.855 63.655 ;
        RECT 137.145 63.485 137.315 63.655 ;
        RECT 137.605 63.485 137.775 63.655 ;
        RECT 138.065 63.485 138.235 63.655 ;
        RECT 138.525 63.485 138.695 63.655 ;
        RECT 138.985 63.485 139.155 63.655 ;
        RECT 50.665 60.765 50.835 60.935 ;
        RECT 51.125 60.765 51.295 60.935 ;
        RECT 51.585 60.765 51.755 60.935 ;
        RECT 52.045 60.765 52.215 60.935 ;
        RECT 52.505 60.765 52.675 60.935 ;
        RECT 52.965 60.765 53.135 60.935 ;
        RECT 53.425 60.765 53.595 60.935 ;
        RECT 53.885 60.765 54.055 60.935 ;
        RECT 54.345 60.765 54.515 60.935 ;
        RECT 54.805 60.765 54.975 60.935 ;
        RECT 55.265 60.765 55.435 60.935 ;
        RECT 55.725 60.765 55.895 60.935 ;
        RECT 56.185 60.765 56.355 60.935 ;
        RECT 56.645 60.765 56.815 60.935 ;
        RECT 57.105 60.765 57.275 60.935 ;
        RECT 57.565 60.765 57.735 60.935 ;
        RECT 58.025 60.765 58.195 60.935 ;
        RECT 58.485 60.765 58.655 60.935 ;
        RECT 58.945 60.765 59.115 60.935 ;
        RECT 59.405 60.765 59.575 60.935 ;
        RECT 59.865 60.765 60.035 60.935 ;
        RECT 60.325 60.765 60.495 60.935 ;
        RECT 60.785 60.765 60.955 60.935 ;
        RECT 61.245 60.765 61.415 60.935 ;
        RECT 61.705 60.765 61.875 60.935 ;
        RECT 62.165 60.765 62.335 60.935 ;
        RECT 62.625 60.765 62.795 60.935 ;
        RECT 63.085 60.765 63.255 60.935 ;
        RECT 63.545 60.765 63.715 60.935 ;
        RECT 64.005 60.765 64.175 60.935 ;
        RECT 64.465 60.765 64.635 60.935 ;
        RECT 64.925 60.765 65.095 60.935 ;
        RECT 65.385 60.765 65.555 60.935 ;
        RECT 65.845 60.765 66.015 60.935 ;
        RECT 66.305 60.765 66.475 60.935 ;
        RECT 66.765 60.765 66.935 60.935 ;
        RECT 67.225 60.765 67.395 60.935 ;
        RECT 67.685 60.765 67.855 60.935 ;
        RECT 68.145 60.765 68.315 60.935 ;
        RECT 68.605 60.765 68.775 60.935 ;
        RECT 69.065 60.765 69.235 60.935 ;
        RECT 69.525 60.765 69.695 60.935 ;
        RECT 69.985 60.765 70.155 60.935 ;
        RECT 70.445 60.765 70.615 60.935 ;
        RECT 70.905 60.765 71.075 60.935 ;
        RECT 71.365 60.765 71.535 60.935 ;
        RECT 71.825 60.765 71.995 60.935 ;
        RECT 72.285 60.765 72.455 60.935 ;
        RECT 72.745 60.765 72.915 60.935 ;
        RECT 73.205 60.765 73.375 60.935 ;
        RECT 73.665 60.765 73.835 60.935 ;
        RECT 74.125 60.765 74.295 60.935 ;
        RECT 74.585 60.765 74.755 60.935 ;
        RECT 75.045 60.765 75.215 60.935 ;
        RECT 75.505 60.765 75.675 60.935 ;
        RECT 75.965 60.765 76.135 60.935 ;
        RECT 76.425 60.765 76.595 60.935 ;
        RECT 76.885 60.765 77.055 60.935 ;
        RECT 77.345 60.765 77.515 60.935 ;
        RECT 77.805 60.765 77.975 60.935 ;
        RECT 78.265 60.765 78.435 60.935 ;
        RECT 78.725 60.765 78.895 60.935 ;
        RECT 79.185 60.765 79.355 60.935 ;
        RECT 79.645 60.765 79.815 60.935 ;
        RECT 80.105 60.765 80.275 60.935 ;
        RECT 80.565 60.765 80.735 60.935 ;
        RECT 81.025 60.765 81.195 60.935 ;
        RECT 81.485 60.765 81.655 60.935 ;
        RECT 81.945 60.765 82.115 60.935 ;
        RECT 82.405 60.765 82.575 60.935 ;
        RECT 82.865 60.765 83.035 60.935 ;
        RECT 83.325 60.765 83.495 60.935 ;
        RECT 83.785 60.765 83.955 60.935 ;
        RECT 84.245 60.765 84.415 60.935 ;
        RECT 84.705 60.765 84.875 60.935 ;
        RECT 85.165 60.765 85.335 60.935 ;
        RECT 85.625 60.765 85.795 60.935 ;
        RECT 86.085 60.765 86.255 60.935 ;
        RECT 86.545 60.765 86.715 60.935 ;
        RECT 87.005 60.765 87.175 60.935 ;
        RECT 87.465 60.765 87.635 60.935 ;
        RECT 87.925 60.765 88.095 60.935 ;
        RECT 88.385 60.765 88.555 60.935 ;
        RECT 88.845 60.765 89.015 60.935 ;
        RECT 89.305 60.765 89.475 60.935 ;
        RECT 89.765 60.765 89.935 60.935 ;
        RECT 90.225 60.765 90.395 60.935 ;
        RECT 90.685 60.765 90.855 60.935 ;
        RECT 91.145 60.765 91.315 60.935 ;
        RECT 91.605 60.765 91.775 60.935 ;
        RECT 92.065 60.765 92.235 60.935 ;
        RECT 92.525 60.765 92.695 60.935 ;
        RECT 92.985 60.765 93.155 60.935 ;
        RECT 93.445 60.765 93.615 60.935 ;
        RECT 93.905 60.765 94.075 60.935 ;
        RECT 94.365 60.765 94.535 60.935 ;
        RECT 94.825 60.765 94.995 60.935 ;
        RECT 95.285 60.765 95.455 60.935 ;
        RECT 95.745 60.765 95.915 60.935 ;
        RECT 96.205 60.765 96.375 60.935 ;
        RECT 96.665 60.765 96.835 60.935 ;
        RECT 97.125 60.765 97.295 60.935 ;
        RECT 97.585 60.765 97.755 60.935 ;
        RECT 98.045 60.765 98.215 60.935 ;
        RECT 98.505 60.765 98.675 60.935 ;
        RECT 98.965 60.765 99.135 60.935 ;
        RECT 99.425 60.765 99.595 60.935 ;
        RECT 99.885 60.765 100.055 60.935 ;
        RECT 100.345 60.765 100.515 60.935 ;
        RECT 100.805 60.765 100.975 60.935 ;
        RECT 101.265 60.765 101.435 60.935 ;
        RECT 101.725 60.765 101.895 60.935 ;
        RECT 102.185 60.765 102.355 60.935 ;
        RECT 102.645 60.765 102.815 60.935 ;
        RECT 103.105 60.765 103.275 60.935 ;
        RECT 103.565 60.765 103.735 60.935 ;
        RECT 104.025 60.765 104.195 60.935 ;
        RECT 104.485 60.765 104.655 60.935 ;
        RECT 104.945 60.765 105.115 60.935 ;
        RECT 105.405 60.765 105.575 60.935 ;
        RECT 105.865 60.765 106.035 60.935 ;
        RECT 106.325 60.765 106.495 60.935 ;
        RECT 106.785 60.765 106.955 60.935 ;
        RECT 107.245 60.765 107.415 60.935 ;
        RECT 107.705 60.765 107.875 60.935 ;
        RECT 108.165 60.765 108.335 60.935 ;
        RECT 108.625 60.765 108.795 60.935 ;
        RECT 109.085 60.765 109.255 60.935 ;
        RECT 109.545 60.765 109.715 60.935 ;
        RECT 110.005 60.765 110.175 60.935 ;
        RECT 110.465 60.765 110.635 60.935 ;
        RECT 110.925 60.765 111.095 60.935 ;
        RECT 111.385 60.765 111.555 60.935 ;
        RECT 111.845 60.765 112.015 60.935 ;
        RECT 112.305 60.765 112.475 60.935 ;
        RECT 112.765 60.765 112.935 60.935 ;
        RECT 113.225 60.765 113.395 60.935 ;
        RECT 113.685 60.765 113.855 60.935 ;
        RECT 114.145 60.765 114.315 60.935 ;
        RECT 114.605 60.765 114.775 60.935 ;
        RECT 115.065 60.765 115.235 60.935 ;
        RECT 115.525 60.765 115.695 60.935 ;
        RECT 115.985 60.765 116.155 60.935 ;
        RECT 116.445 60.765 116.615 60.935 ;
        RECT 116.905 60.765 117.075 60.935 ;
        RECT 117.365 60.765 117.535 60.935 ;
        RECT 117.825 60.765 117.995 60.935 ;
        RECT 118.285 60.765 118.455 60.935 ;
        RECT 118.745 60.765 118.915 60.935 ;
        RECT 119.205 60.765 119.375 60.935 ;
        RECT 119.665 60.765 119.835 60.935 ;
        RECT 120.125 60.765 120.295 60.935 ;
        RECT 120.585 60.765 120.755 60.935 ;
        RECT 121.045 60.765 121.215 60.935 ;
        RECT 121.505 60.765 121.675 60.935 ;
        RECT 121.965 60.765 122.135 60.935 ;
        RECT 122.425 60.765 122.595 60.935 ;
        RECT 122.885 60.765 123.055 60.935 ;
        RECT 123.345 60.765 123.515 60.935 ;
        RECT 123.805 60.765 123.975 60.935 ;
        RECT 124.265 60.765 124.435 60.935 ;
        RECT 124.725 60.765 124.895 60.935 ;
        RECT 125.185 60.765 125.355 60.935 ;
        RECT 125.645 60.765 125.815 60.935 ;
        RECT 126.105 60.765 126.275 60.935 ;
        RECT 126.565 60.765 126.735 60.935 ;
        RECT 127.025 60.765 127.195 60.935 ;
        RECT 127.485 60.765 127.655 60.935 ;
        RECT 127.945 60.765 128.115 60.935 ;
        RECT 128.405 60.765 128.575 60.935 ;
        RECT 128.865 60.765 129.035 60.935 ;
        RECT 129.325 60.765 129.495 60.935 ;
        RECT 129.785 60.765 129.955 60.935 ;
        RECT 130.245 60.765 130.415 60.935 ;
        RECT 130.705 60.765 130.875 60.935 ;
        RECT 131.165 60.765 131.335 60.935 ;
        RECT 131.625 60.765 131.795 60.935 ;
        RECT 132.085 60.765 132.255 60.935 ;
        RECT 132.545 60.765 132.715 60.935 ;
        RECT 133.005 60.765 133.175 60.935 ;
        RECT 133.465 60.765 133.635 60.935 ;
        RECT 133.925 60.765 134.095 60.935 ;
        RECT 134.385 60.765 134.555 60.935 ;
        RECT 134.845 60.765 135.015 60.935 ;
        RECT 135.305 60.765 135.475 60.935 ;
        RECT 135.765 60.765 135.935 60.935 ;
        RECT 136.225 60.765 136.395 60.935 ;
        RECT 136.685 60.765 136.855 60.935 ;
        RECT 137.145 60.765 137.315 60.935 ;
        RECT 137.605 60.765 137.775 60.935 ;
        RECT 138.065 60.765 138.235 60.935 ;
        RECT 138.525 60.765 138.695 60.935 ;
        RECT 138.985 60.765 139.155 60.935 ;
      LAYER met1 ;
        RECT 50.520 136.770 140.095 137.250 ;
        RECT 50.520 134.050 139.300 134.530 ;
        RECT 50.520 131.330 140.095 131.810 ;
        RECT 50.520 128.610 139.300 129.090 ;
        RECT 50.520 125.890 140.095 126.370 ;
        RECT 50.520 123.170 139.300 123.650 ;
        RECT 50.520 120.450 140.095 120.930 ;
        RECT 50.520 117.730 139.300 118.210 ;
        RECT 50.520 115.010 140.095 115.490 ;
        RECT 50.520 112.290 139.300 112.770 ;
        RECT 50.520 109.570 140.095 110.050 ;
        RECT 63.930 108.690 64.250 108.750 ;
        RECT 65.325 108.690 65.615 108.735 ;
        RECT 63.930 108.550 65.615 108.690 ;
        RECT 63.930 108.490 64.250 108.550 ;
        RECT 65.325 108.505 65.615 108.550 ;
        RECT 65.785 108.690 66.075 108.735 ;
        RECT 66.705 108.690 66.995 108.735 ;
        RECT 65.785 108.550 66.995 108.690 ;
        RECT 65.785 108.505 66.075 108.550 ;
        RECT 66.705 108.505 66.995 108.550 ;
        RECT 50.520 106.850 139.300 107.330 ;
        RECT 57.965 105.970 58.255 106.015 ;
        RECT 61.185 105.970 61.475 106.015 ;
        RECT 57.965 105.830 61.475 105.970 ;
        RECT 57.965 105.785 58.255 105.830 ;
        RECT 61.185 105.785 61.475 105.830 ;
        RECT 57.030 105.630 57.350 105.690 ;
        RECT 57.505 105.630 57.795 105.675 ;
        RECT 57.030 105.490 57.795 105.630 ;
        RECT 57.030 105.430 57.350 105.490 ;
        RECT 57.505 105.445 57.795 105.490 ;
        RECT 58.425 105.630 58.715 105.675 ;
        RECT 60.250 105.630 60.570 105.690 ;
        RECT 58.425 105.490 60.570 105.630 ;
        RECT 58.425 105.445 58.715 105.490 ;
        RECT 60.250 105.430 60.570 105.490 ;
        RECT 62.105 105.630 62.395 105.675 ;
        RECT 62.550 105.630 62.870 105.690 ;
        RECT 62.105 105.490 62.870 105.630 ;
        RECT 62.105 105.445 62.395 105.490 ;
        RECT 62.550 105.430 62.870 105.490 ;
        RECT 58.870 105.090 59.190 105.350 ;
        RECT 50.520 104.130 140.095 104.610 ;
        RECT 52.905 103.930 53.195 103.975 ;
        RECT 57.030 103.930 57.350 103.990 ;
        RECT 52.905 103.790 57.350 103.930 ;
        RECT 52.905 103.745 53.195 103.790 ;
        RECT 57.030 103.730 57.350 103.790 ;
        RECT 48.750 103.250 49.070 103.310 ;
        RECT 51.985 103.250 52.275 103.295 ;
        RECT 48.750 103.110 52.275 103.250 ;
        RECT 57.120 103.250 57.260 103.730 ;
        RECT 61.645 103.590 61.935 103.635 ;
        RECT 63.025 103.590 63.315 103.635 ;
        RECT 63.470 103.590 63.790 103.650 ;
        RECT 61.645 103.450 63.790 103.590 ;
        RECT 61.645 103.405 61.935 103.450 ;
        RECT 63.025 103.405 63.315 103.450 ;
        RECT 63.470 103.390 63.790 103.450 ;
        RECT 59.805 103.250 60.095 103.295 ;
        RECT 57.120 103.110 60.095 103.250 ;
        RECT 48.750 103.050 49.070 103.110 ;
        RECT 51.985 103.065 52.275 103.110 ;
        RECT 59.805 103.065 60.095 103.110 ;
        RECT 60.250 103.250 60.570 103.310 ;
        RECT 61.185 103.250 61.475 103.295 ;
        RECT 60.250 103.110 61.475 103.250 ;
        RECT 60.250 103.050 60.570 103.110 ;
        RECT 61.185 103.065 61.475 103.110 ;
        RECT 62.105 103.250 62.400 103.295 ;
        RECT 65.340 103.250 65.630 103.295 ;
        RECT 62.105 103.110 65.630 103.250 ;
        RECT 62.105 103.065 62.400 103.110 ;
        RECT 65.340 103.065 65.630 103.110 ;
        RECT 61.260 102.570 61.400 103.065 ;
        RECT 62.550 102.710 62.870 102.970 ;
        RECT 63.930 102.710 64.250 102.970 ;
        RECT 64.020 102.570 64.160 102.710 ;
        RECT 61.260 102.430 64.160 102.570 ;
        RECT 50.520 101.410 139.300 101.890 ;
        RECT 51.985 100.190 52.275 100.235 ;
        RECT 58.870 100.190 59.190 100.250 ;
        RECT 51.985 100.050 59.190 100.190 ;
        RECT 51.985 100.005 52.275 100.050 ;
        RECT 58.870 99.990 59.190 100.050 ;
        RECT 52.905 99.510 53.195 99.555 ;
        RECT 58.410 99.510 58.730 99.570 ;
        RECT 52.905 99.370 58.730 99.510 ;
        RECT 52.905 99.325 53.195 99.370 ;
        RECT 58.410 99.310 58.730 99.370 ;
        RECT 50.520 98.690 140.095 99.170 ;
        RECT 61.645 98.490 61.935 98.535 ;
        RECT 62.550 98.490 62.870 98.550 ;
        RECT 61.645 98.350 62.870 98.490 ;
        RECT 61.645 98.305 61.935 98.350 ;
        RECT 62.550 98.290 62.870 98.350 ;
        RECT 60.250 97.810 60.570 97.870 ;
        RECT 60.725 97.810 61.015 97.855 ;
        RECT 60.250 97.670 61.015 97.810 ;
        RECT 60.250 97.610 60.570 97.670 ;
        RECT 60.725 97.625 61.015 97.670 ;
        RECT 50.520 95.970 139.300 96.450 ;
        RECT 58.410 94.750 58.730 94.810 ;
        RECT 61.645 94.750 61.935 94.795 ;
        RECT 58.410 94.610 61.935 94.750 ;
        RECT 58.410 94.550 58.730 94.610 ;
        RECT 61.645 94.565 61.935 94.610 ;
        RECT 62.565 94.750 62.855 94.795 ;
        RECT 63.930 94.750 64.250 94.810 ;
        RECT 62.565 94.610 64.250 94.750 ;
        RECT 62.565 94.565 62.855 94.610 ;
        RECT 63.930 94.550 64.250 94.610 ;
        RECT 57.950 94.070 58.270 94.130 ;
        RECT 61.645 94.070 61.935 94.115 ;
        RECT 66.230 94.070 66.550 94.130 ;
        RECT 57.950 93.930 66.550 94.070 ;
        RECT 57.950 93.870 58.270 93.930 ;
        RECT 61.645 93.885 61.935 93.930 ;
        RECT 66.230 93.870 66.550 93.930 ;
        RECT 50.520 93.250 140.095 93.730 ;
        RECT 57.950 92.850 58.270 93.110 ;
        RECT 58.410 92.850 58.730 93.110 ;
        RECT 60.250 93.050 60.570 93.110 ;
        RECT 60.725 93.050 61.015 93.095 ;
        RECT 60.250 92.910 61.015 93.050 ;
        RECT 60.250 92.850 60.570 92.910 ;
        RECT 60.725 92.865 61.015 92.910 ;
        RECT 63.025 92.710 63.315 92.755 ;
        RECT 66.705 92.710 66.995 92.755 ;
        RECT 63.025 92.570 66.995 92.710 ;
        RECT 63.025 92.525 63.315 92.570 ;
        RECT 66.705 92.525 66.995 92.570 ;
        RECT 62.550 92.170 62.870 92.430 ;
        RECT 64.865 92.370 65.155 92.415 ;
        RECT 63.560 92.230 65.155 92.370 ;
        RECT 63.560 92.090 63.700 92.230 ;
        RECT 64.865 92.185 65.155 92.230 ;
        RECT 66.230 92.170 66.550 92.430 ;
        RECT 57.505 92.030 57.795 92.075 ;
        RECT 63.470 92.030 63.790 92.090 ;
        RECT 57.505 91.890 63.790 92.030 ;
        RECT 57.505 91.845 57.795 91.890 ;
        RECT 63.470 91.830 63.790 91.890 ;
        RECT 60.250 91.150 60.570 91.410 ;
        RECT 50.520 90.530 139.300 91.010 ;
        RECT 62.105 90.330 62.395 90.375 ;
        RECT 62.550 90.330 62.870 90.390 ;
        RECT 62.105 90.190 62.870 90.330 ;
        RECT 62.105 90.145 62.395 90.190 ;
        RECT 62.550 90.130 62.870 90.190 ;
        RECT 58.870 89.650 59.190 89.710 ;
        RECT 58.870 89.510 61.860 89.650 ;
        RECT 58.870 89.450 59.190 89.510 ;
        RECT 60.250 89.110 60.570 89.370 ;
        RECT 61.720 89.355 61.860 89.510 ;
        RECT 61.645 89.125 61.935 89.355 ;
        RECT 50.520 87.810 140.095 88.290 ;
        RECT 50.520 85.090 139.300 85.570 ;
        RECT 50.520 82.370 140.095 82.850 ;
        RECT 50.520 79.650 139.300 80.130 ;
        RECT 50.520 76.930 140.095 77.410 ;
        RECT 50.520 74.210 139.300 74.690 ;
        RECT 50.520 71.490 140.095 71.970 ;
        RECT 50.520 68.770 139.300 69.250 ;
        RECT 50.520 66.050 140.095 66.530 ;
        RECT 50.520 63.330 139.300 63.810 ;
        RECT 50.520 60.610 140.095 61.090 ;
      LAYER via ;
        RECT 71.940 136.880 72.200 137.140 ;
        RECT 72.260 136.880 72.520 137.140 ;
        RECT 72.580 136.880 72.840 137.140 ;
        RECT 72.900 136.880 73.160 137.140 ;
        RECT 73.220 136.880 73.480 137.140 ;
        RECT 94.135 136.880 94.395 137.140 ;
        RECT 94.455 136.880 94.715 137.140 ;
        RECT 94.775 136.880 95.035 137.140 ;
        RECT 95.095 136.880 95.355 137.140 ;
        RECT 95.415 136.880 95.675 137.140 ;
        RECT 116.330 136.880 116.590 137.140 ;
        RECT 116.650 136.880 116.910 137.140 ;
        RECT 116.970 136.880 117.230 137.140 ;
        RECT 117.290 136.880 117.550 137.140 ;
        RECT 117.610 136.880 117.870 137.140 ;
        RECT 138.525 136.880 138.785 137.140 ;
        RECT 138.845 136.880 139.105 137.140 ;
        RECT 139.165 136.880 139.425 137.140 ;
        RECT 139.485 136.880 139.745 137.140 ;
        RECT 139.805 136.880 140.065 137.140 ;
        RECT 60.845 134.160 61.105 134.420 ;
        RECT 61.165 134.160 61.425 134.420 ;
        RECT 61.485 134.160 61.745 134.420 ;
        RECT 61.805 134.160 62.065 134.420 ;
        RECT 62.125 134.160 62.385 134.420 ;
        RECT 83.040 134.160 83.300 134.420 ;
        RECT 83.360 134.160 83.620 134.420 ;
        RECT 83.680 134.160 83.940 134.420 ;
        RECT 84.000 134.160 84.260 134.420 ;
        RECT 84.320 134.160 84.580 134.420 ;
        RECT 105.235 134.160 105.495 134.420 ;
        RECT 105.555 134.160 105.815 134.420 ;
        RECT 105.875 134.160 106.135 134.420 ;
        RECT 106.195 134.160 106.455 134.420 ;
        RECT 106.515 134.160 106.775 134.420 ;
        RECT 127.430 134.160 127.690 134.420 ;
        RECT 127.750 134.160 128.010 134.420 ;
        RECT 128.070 134.160 128.330 134.420 ;
        RECT 128.390 134.160 128.650 134.420 ;
        RECT 128.710 134.160 128.970 134.420 ;
        RECT 71.940 131.440 72.200 131.700 ;
        RECT 72.260 131.440 72.520 131.700 ;
        RECT 72.580 131.440 72.840 131.700 ;
        RECT 72.900 131.440 73.160 131.700 ;
        RECT 73.220 131.440 73.480 131.700 ;
        RECT 94.135 131.440 94.395 131.700 ;
        RECT 94.455 131.440 94.715 131.700 ;
        RECT 94.775 131.440 95.035 131.700 ;
        RECT 95.095 131.440 95.355 131.700 ;
        RECT 95.415 131.440 95.675 131.700 ;
        RECT 116.330 131.440 116.590 131.700 ;
        RECT 116.650 131.440 116.910 131.700 ;
        RECT 116.970 131.440 117.230 131.700 ;
        RECT 117.290 131.440 117.550 131.700 ;
        RECT 117.610 131.440 117.870 131.700 ;
        RECT 138.525 131.440 138.785 131.700 ;
        RECT 138.845 131.440 139.105 131.700 ;
        RECT 139.165 131.440 139.425 131.700 ;
        RECT 139.485 131.440 139.745 131.700 ;
        RECT 139.805 131.440 140.065 131.700 ;
        RECT 60.845 128.720 61.105 128.980 ;
        RECT 61.165 128.720 61.425 128.980 ;
        RECT 61.485 128.720 61.745 128.980 ;
        RECT 61.805 128.720 62.065 128.980 ;
        RECT 62.125 128.720 62.385 128.980 ;
        RECT 83.040 128.720 83.300 128.980 ;
        RECT 83.360 128.720 83.620 128.980 ;
        RECT 83.680 128.720 83.940 128.980 ;
        RECT 84.000 128.720 84.260 128.980 ;
        RECT 84.320 128.720 84.580 128.980 ;
        RECT 105.235 128.720 105.495 128.980 ;
        RECT 105.555 128.720 105.815 128.980 ;
        RECT 105.875 128.720 106.135 128.980 ;
        RECT 106.195 128.720 106.455 128.980 ;
        RECT 106.515 128.720 106.775 128.980 ;
        RECT 127.430 128.720 127.690 128.980 ;
        RECT 127.750 128.720 128.010 128.980 ;
        RECT 128.070 128.720 128.330 128.980 ;
        RECT 128.390 128.720 128.650 128.980 ;
        RECT 128.710 128.720 128.970 128.980 ;
        RECT 71.940 126.000 72.200 126.260 ;
        RECT 72.260 126.000 72.520 126.260 ;
        RECT 72.580 126.000 72.840 126.260 ;
        RECT 72.900 126.000 73.160 126.260 ;
        RECT 73.220 126.000 73.480 126.260 ;
        RECT 94.135 126.000 94.395 126.260 ;
        RECT 94.455 126.000 94.715 126.260 ;
        RECT 94.775 126.000 95.035 126.260 ;
        RECT 95.095 126.000 95.355 126.260 ;
        RECT 95.415 126.000 95.675 126.260 ;
        RECT 116.330 126.000 116.590 126.260 ;
        RECT 116.650 126.000 116.910 126.260 ;
        RECT 116.970 126.000 117.230 126.260 ;
        RECT 117.290 126.000 117.550 126.260 ;
        RECT 117.610 126.000 117.870 126.260 ;
        RECT 138.525 126.000 138.785 126.260 ;
        RECT 138.845 126.000 139.105 126.260 ;
        RECT 139.165 126.000 139.425 126.260 ;
        RECT 139.485 126.000 139.745 126.260 ;
        RECT 139.805 126.000 140.065 126.260 ;
        RECT 60.845 123.280 61.105 123.540 ;
        RECT 61.165 123.280 61.425 123.540 ;
        RECT 61.485 123.280 61.745 123.540 ;
        RECT 61.805 123.280 62.065 123.540 ;
        RECT 62.125 123.280 62.385 123.540 ;
        RECT 83.040 123.280 83.300 123.540 ;
        RECT 83.360 123.280 83.620 123.540 ;
        RECT 83.680 123.280 83.940 123.540 ;
        RECT 84.000 123.280 84.260 123.540 ;
        RECT 84.320 123.280 84.580 123.540 ;
        RECT 105.235 123.280 105.495 123.540 ;
        RECT 105.555 123.280 105.815 123.540 ;
        RECT 105.875 123.280 106.135 123.540 ;
        RECT 106.195 123.280 106.455 123.540 ;
        RECT 106.515 123.280 106.775 123.540 ;
        RECT 127.430 123.280 127.690 123.540 ;
        RECT 127.750 123.280 128.010 123.540 ;
        RECT 128.070 123.280 128.330 123.540 ;
        RECT 128.390 123.280 128.650 123.540 ;
        RECT 128.710 123.280 128.970 123.540 ;
        RECT 71.940 120.560 72.200 120.820 ;
        RECT 72.260 120.560 72.520 120.820 ;
        RECT 72.580 120.560 72.840 120.820 ;
        RECT 72.900 120.560 73.160 120.820 ;
        RECT 73.220 120.560 73.480 120.820 ;
        RECT 94.135 120.560 94.395 120.820 ;
        RECT 94.455 120.560 94.715 120.820 ;
        RECT 94.775 120.560 95.035 120.820 ;
        RECT 95.095 120.560 95.355 120.820 ;
        RECT 95.415 120.560 95.675 120.820 ;
        RECT 116.330 120.560 116.590 120.820 ;
        RECT 116.650 120.560 116.910 120.820 ;
        RECT 116.970 120.560 117.230 120.820 ;
        RECT 117.290 120.560 117.550 120.820 ;
        RECT 117.610 120.560 117.870 120.820 ;
        RECT 138.525 120.560 138.785 120.820 ;
        RECT 138.845 120.560 139.105 120.820 ;
        RECT 139.165 120.560 139.425 120.820 ;
        RECT 139.485 120.560 139.745 120.820 ;
        RECT 139.805 120.560 140.065 120.820 ;
        RECT 60.845 117.840 61.105 118.100 ;
        RECT 61.165 117.840 61.425 118.100 ;
        RECT 61.485 117.840 61.745 118.100 ;
        RECT 61.805 117.840 62.065 118.100 ;
        RECT 62.125 117.840 62.385 118.100 ;
        RECT 83.040 117.840 83.300 118.100 ;
        RECT 83.360 117.840 83.620 118.100 ;
        RECT 83.680 117.840 83.940 118.100 ;
        RECT 84.000 117.840 84.260 118.100 ;
        RECT 84.320 117.840 84.580 118.100 ;
        RECT 105.235 117.840 105.495 118.100 ;
        RECT 105.555 117.840 105.815 118.100 ;
        RECT 105.875 117.840 106.135 118.100 ;
        RECT 106.195 117.840 106.455 118.100 ;
        RECT 106.515 117.840 106.775 118.100 ;
        RECT 127.430 117.840 127.690 118.100 ;
        RECT 127.750 117.840 128.010 118.100 ;
        RECT 128.070 117.840 128.330 118.100 ;
        RECT 128.390 117.840 128.650 118.100 ;
        RECT 128.710 117.840 128.970 118.100 ;
        RECT 71.940 115.120 72.200 115.380 ;
        RECT 72.260 115.120 72.520 115.380 ;
        RECT 72.580 115.120 72.840 115.380 ;
        RECT 72.900 115.120 73.160 115.380 ;
        RECT 73.220 115.120 73.480 115.380 ;
        RECT 94.135 115.120 94.395 115.380 ;
        RECT 94.455 115.120 94.715 115.380 ;
        RECT 94.775 115.120 95.035 115.380 ;
        RECT 95.095 115.120 95.355 115.380 ;
        RECT 95.415 115.120 95.675 115.380 ;
        RECT 116.330 115.120 116.590 115.380 ;
        RECT 116.650 115.120 116.910 115.380 ;
        RECT 116.970 115.120 117.230 115.380 ;
        RECT 117.290 115.120 117.550 115.380 ;
        RECT 117.610 115.120 117.870 115.380 ;
        RECT 138.525 115.120 138.785 115.380 ;
        RECT 138.845 115.120 139.105 115.380 ;
        RECT 139.165 115.120 139.425 115.380 ;
        RECT 139.485 115.120 139.745 115.380 ;
        RECT 139.805 115.120 140.065 115.380 ;
        RECT 60.845 112.400 61.105 112.660 ;
        RECT 61.165 112.400 61.425 112.660 ;
        RECT 61.485 112.400 61.745 112.660 ;
        RECT 61.805 112.400 62.065 112.660 ;
        RECT 62.125 112.400 62.385 112.660 ;
        RECT 83.040 112.400 83.300 112.660 ;
        RECT 83.360 112.400 83.620 112.660 ;
        RECT 83.680 112.400 83.940 112.660 ;
        RECT 84.000 112.400 84.260 112.660 ;
        RECT 84.320 112.400 84.580 112.660 ;
        RECT 105.235 112.400 105.495 112.660 ;
        RECT 105.555 112.400 105.815 112.660 ;
        RECT 105.875 112.400 106.135 112.660 ;
        RECT 106.195 112.400 106.455 112.660 ;
        RECT 106.515 112.400 106.775 112.660 ;
        RECT 127.430 112.400 127.690 112.660 ;
        RECT 127.750 112.400 128.010 112.660 ;
        RECT 128.070 112.400 128.330 112.660 ;
        RECT 128.390 112.400 128.650 112.660 ;
        RECT 128.710 112.400 128.970 112.660 ;
        RECT 71.940 109.680 72.200 109.940 ;
        RECT 72.260 109.680 72.520 109.940 ;
        RECT 72.580 109.680 72.840 109.940 ;
        RECT 72.900 109.680 73.160 109.940 ;
        RECT 73.220 109.680 73.480 109.940 ;
        RECT 94.135 109.680 94.395 109.940 ;
        RECT 94.455 109.680 94.715 109.940 ;
        RECT 94.775 109.680 95.035 109.940 ;
        RECT 95.095 109.680 95.355 109.940 ;
        RECT 95.415 109.680 95.675 109.940 ;
        RECT 116.330 109.680 116.590 109.940 ;
        RECT 116.650 109.680 116.910 109.940 ;
        RECT 116.970 109.680 117.230 109.940 ;
        RECT 117.290 109.680 117.550 109.940 ;
        RECT 117.610 109.680 117.870 109.940 ;
        RECT 138.525 109.680 138.785 109.940 ;
        RECT 138.845 109.680 139.105 109.940 ;
        RECT 139.165 109.680 139.425 109.940 ;
        RECT 139.485 109.680 139.745 109.940 ;
        RECT 139.805 109.680 140.065 109.940 ;
        RECT 63.960 108.490 64.220 108.750 ;
        RECT 60.845 106.960 61.105 107.220 ;
        RECT 61.165 106.960 61.425 107.220 ;
        RECT 61.485 106.960 61.745 107.220 ;
        RECT 61.805 106.960 62.065 107.220 ;
        RECT 62.125 106.960 62.385 107.220 ;
        RECT 83.040 106.960 83.300 107.220 ;
        RECT 83.360 106.960 83.620 107.220 ;
        RECT 83.680 106.960 83.940 107.220 ;
        RECT 84.000 106.960 84.260 107.220 ;
        RECT 84.320 106.960 84.580 107.220 ;
        RECT 105.235 106.960 105.495 107.220 ;
        RECT 105.555 106.960 105.815 107.220 ;
        RECT 105.875 106.960 106.135 107.220 ;
        RECT 106.195 106.960 106.455 107.220 ;
        RECT 106.515 106.960 106.775 107.220 ;
        RECT 127.430 106.960 127.690 107.220 ;
        RECT 127.750 106.960 128.010 107.220 ;
        RECT 128.070 106.960 128.330 107.220 ;
        RECT 128.390 106.960 128.650 107.220 ;
        RECT 128.710 106.960 128.970 107.220 ;
        RECT 57.060 105.430 57.320 105.690 ;
        RECT 60.280 105.430 60.540 105.690 ;
        RECT 62.580 105.430 62.840 105.690 ;
        RECT 58.900 105.090 59.160 105.350 ;
        RECT 71.940 104.240 72.200 104.500 ;
        RECT 72.260 104.240 72.520 104.500 ;
        RECT 72.580 104.240 72.840 104.500 ;
        RECT 72.900 104.240 73.160 104.500 ;
        RECT 73.220 104.240 73.480 104.500 ;
        RECT 94.135 104.240 94.395 104.500 ;
        RECT 94.455 104.240 94.715 104.500 ;
        RECT 94.775 104.240 95.035 104.500 ;
        RECT 95.095 104.240 95.355 104.500 ;
        RECT 95.415 104.240 95.675 104.500 ;
        RECT 116.330 104.240 116.590 104.500 ;
        RECT 116.650 104.240 116.910 104.500 ;
        RECT 116.970 104.240 117.230 104.500 ;
        RECT 117.290 104.240 117.550 104.500 ;
        RECT 117.610 104.240 117.870 104.500 ;
        RECT 138.525 104.240 138.785 104.500 ;
        RECT 138.845 104.240 139.105 104.500 ;
        RECT 139.165 104.240 139.425 104.500 ;
        RECT 139.485 104.240 139.745 104.500 ;
        RECT 139.805 104.240 140.065 104.500 ;
        RECT 57.060 103.730 57.320 103.990 ;
        RECT 48.780 103.050 49.040 103.310 ;
        RECT 63.500 103.390 63.760 103.650 ;
        RECT 60.280 103.050 60.540 103.310 ;
        RECT 62.580 102.710 62.840 102.970 ;
        RECT 63.960 102.710 64.220 102.970 ;
        RECT 60.845 101.520 61.105 101.780 ;
        RECT 61.165 101.520 61.425 101.780 ;
        RECT 61.485 101.520 61.745 101.780 ;
        RECT 61.805 101.520 62.065 101.780 ;
        RECT 62.125 101.520 62.385 101.780 ;
        RECT 83.040 101.520 83.300 101.780 ;
        RECT 83.360 101.520 83.620 101.780 ;
        RECT 83.680 101.520 83.940 101.780 ;
        RECT 84.000 101.520 84.260 101.780 ;
        RECT 84.320 101.520 84.580 101.780 ;
        RECT 105.235 101.520 105.495 101.780 ;
        RECT 105.555 101.520 105.815 101.780 ;
        RECT 105.875 101.520 106.135 101.780 ;
        RECT 106.195 101.520 106.455 101.780 ;
        RECT 106.515 101.520 106.775 101.780 ;
        RECT 127.430 101.520 127.690 101.780 ;
        RECT 127.750 101.520 128.010 101.780 ;
        RECT 128.070 101.520 128.330 101.780 ;
        RECT 128.390 101.520 128.650 101.780 ;
        RECT 128.710 101.520 128.970 101.780 ;
        RECT 58.900 99.990 59.160 100.250 ;
        RECT 58.440 99.310 58.700 99.570 ;
        RECT 71.940 98.800 72.200 99.060 ;
        RECT 72.260 98.800 72.520 99.060 ;
        RECT 72.580 98.800 72.840 99.060 ;
        RECT 72.900 98.800 73.160 99.060 ;
        RECT 73.220 98.800 73.480 99.060 ;
        RECT 94.135 98.800 94.395 99.060 ;
        RECT 94.455 98.800 94.715 99.060 ;
        RECT 94.775 98.800 95.035 99.060 ;
        RECT 95.095 98.800 95.355 99.060 ;
        RECT 95.415 98.800 95.675 99.060 ;
        RECT 116.330 98.800 116.590 99.060 ;
        RECT 116.650 98.800 116.910 99.060 ;
        RECT 116.970 98.800 117.230 99.060 ;
        RECT 117.290 98.800 117.550 99.060 ;
        RECT 117.610 98.800 117.870 99.060 ;
        RECT 138.525 98.800 138.785 99.060 ;
        RECT 138.845 98.800 139.105 99.060 ;
        RECT 139.165 98.800 139.425 99.060 ;
        RECT 139.485 98.800 139.745 99.060 ;
        RECT 139.805 98.800 140.065 99.060 ;
        RECT 62.580 98.290 62.840 98.550 ;
        RECT 60.280 97.610 60.540 97.870 ;
        RECT 60.845 96.080 61.105 96.340 ;
        RECT 61.165 96.080 61.425 96.340 ;
        RECT 61.485 96.080 61.745 96.340 ;
        RECT 61.805 96.080 62.065 96.340 ;
        RECT 62.125 96.080 62.385 96.340 ;
        RECT 83.040 96.080 83.300 96.340 ;
        RECT 83.360 96.080 83.620 96.340 ;
        RECT 83.680 96.080 83.940 96.340 ;
        RECT 84.000 96.080 84.260 96.340 ;
        RECT 84.320 96.080 84.580 96.340 ;
        RECT 105.235 96.080 105.495 96.340 ;
        RECT 105.555 96.080 105.815 96.340 ;
        RECT 105.875 96.080 106.135 96.340 ;
        RECT 106.195 96.080 106.455 96.340 ;
        RECT 106.515 96.080 106.775 96.340 ;
        RECT 127.430 96.080 127.690 96.340 ;
        RECT 127.750 96.080 128.010 96.340 ;
        RECT 128.070 96.080 128.330 96.340 ;
        RECT 128.390 96.080 128.650 96.340 ;
        RECT 128.710 96.080 128.970 96.340 ;
        RECT 58.440 94.550 58.700 94.810 ;
        RECT 63.960 94.550 64.220 94.810 ;
        RECT 57.980 93.870 58.240 94.130 ;
        RECT 66.260 93.870 66.520 94.130 ;
        RECT 71.940 93.360 72.200 93.620 ;
        RECT 72.260 93.360 72.520 93.620 ;
        RECT 72.580 93.360 72.840 93.620 ;
        RECT 72.900 93.360 73.160 93.620 ;
        RECT 73.220 93.360 73.480 93.620 ;
        RECT 94.135 93.360 94.395 93.620 ;
        RECT 94.455 93.360 94.715 93.620 ;
        RECT 94.775 93.360 95.035 93.620 ;
        RECT 95.095 93.360 95.355 93.620 ;
        RECT 95.415 93.360 95.675 93.620 ;
        RECT 116.330 93.360 116.590 93.620 ;
        RECT 116.650 93.360 116.910 93.620 ;
        RECT 116.970 93.360 117.230 93.620 ;
        RECT 117.290 93.360 117.550 93.620 ;
        RECT 117.610 93.360 117.870 93.620 ;
        RECT 138.525 93.360 138.785 93.620 ;
        RECT 138.845 93.360 139.105 93.620 ;
        RECT 139.165 93.360 139.425 93.620 ;
        RECT 139.485 93.360 139.745 93.620 ;
        RECT 139.805 93.360 140.065 93.620 ;
        RECT 57.980 92.850 58.240 93.110 ;
        RECT 58.440 92.850 58.700 93.110 ;
        RECT 60.280 92.850 60.540 93.110 ;
        RECT 62.580 92.170 62.840 92.430 ;
        RECT 66.260 92.170 66.520 92.430 ;
        RECT 63.500 91.830 63.760 92.090 ;
        RECT 60.280 91.150 60.540 91.410 ;
        RECT 60.845 90.640 61.105 90.900 ;
        RECT 61.165 90.640 61.425 90.900 ;
        RECT 61.485 90.640 61.745 90.900 ;
        RECT 61.805 90.640 62.065 90.900 ;
        RECT 62.125 90.640 62.385 90.900 ;
        RECT 83.040 90.640 83.300 90.900 ;
        RECT 83.360 90.640 83.620 90.900 ;
        RECT 83.680 90.640 83.940 90.900 ;
        RECT 84.000 90.640 84.260 90.900 ;
        RECT 84.320 90.640 84.580 90.900 ;
        RECT 105.235 90.640 105.495 90.900 ;
        RECT 105.555 90.640 105.815 90.900 ;
        RECT 105.875 90.640 106.135 90.900 ;
        RECT 106.195 90.640 106.455 90.900 ;
        RECT 106.515 90.640 106.775 90.900 ;
        RECT 127.430 90.640 127.690 90.900 ;
        RECT 127.750 90.640 128.010 90.900 ;
        RECT 128.070 90.640 128.330 90.900 ;
        RECT 128.390 90.640 128.650 90.900 ;
        RECT 128.710 90.640 128.970 90.900 ;
        RECT 62.580 90.130 62.840 90.390 ;
        RECT 58.900 89.450 59.160 89.710 ;
        RECT 60.280 89.110 60.540 89.370 ;
        RECT 71.940 87.920 72.200 88.180 ;
        RECT 72.260 87.920 72.520 88.180 ;
        RECT 72.580 87.920 72.840 88.180 ;
        RECT 72.900 87.920 73.160 88.180 ;
        RECT 73.220 87.920 73.480 88.180 ;
        RECT 94.135 87.920 94.395 88.180 ;
        RECT 94.455 87.920 94.715 88.180 ;
        RECT 94.775 87.920 95.035 88.180 ;
        RECT 95.095 87.920 95.355 88.180 ;
        RECT 95.415 87.920 95.675 88.180 ;
        RECT 116.330 87.920 116.590 88.180 ;
        RECT 116.650 87.920 116.910 88.180 ;
        RECT 116.970 87.920 117.230 88.180 ;
        RECT 117.290 87.920 117.550 88.180 ;
        RECT 117.610 87.920 117.870 88.180 ;
        RECT 138.525 87.920 138.785 88.180 ;
        RECT 138.845 87.920 139.105 88.180 ;
        RECT 139.165 87.920 139.425 88.180 ;
        RECT 139.485 87.920 139.745 88.180 ;
        RECT 139.805 87.920 140.065 88.180 ;
        RECT 60.845 85.200 61.105 85.460 ;
        RECT 61.165 85.200 61.425 85.460 ;
        RECT 61.485 85.200 61.745 85.460 ;
        RECT 61.805 85.200 62.065 85.460 ;
        RECT 62.125 85.200 62.385 85.460 ;
        RECT 83.040 85.200 83.300 85.460 ;
        RECT 83.360 85.200 83.620 85.460 ;
        RECT 83.680 85.200 83.940 85.460 ;
        RECT 84.000 85.200 84.260 85.460 ;
        RECT 84.320 85.200 84.580 85.460 ;
        RECT 105.235 85.200 105.495 85.460 ;
        RECT 105.555 85.200 105.815 85.460 ;
        RECT 105.875 85.200 106.135 85.460 ;
        RECT 106.195 85.200 106.455 85.460 ;
        RECT 106.515 85.200 106.775 85.460 ;
        RECT 127.430 85.200 127.690 85.460 ;
        RECT 127.750 85.200 128.010 85.460 ;
        RECT 128.070 85.200 128.330 85.460 ;
        RECT 128.390 85.200 128.650 85.460 ;
        RECT 128.710 85.200 128.970 85.460 ;
        RECT 71.940 82.480 72.200 82.740 ;
        RECT 72.260 82.480 72.520 82.740 ;
        RECT 72.580 82.480 72.840 82.740 ;
        RECT 72.900 82.480 73.160 82.740 ;
        RECT 73.220 82.480 73.480 82.740 ;
        RECT 94.135 82.480 94.395 82.740 ;
        RECT 94.455 82.480 94.715 82.740 ;
        RECT 94.775 82.480 95.035 82.740 ;
        RECT 95.095 82.480 95.355 82.740 ;
        RECT 95.415 82.480 95.675 82.740 ;
        RECT 116.330 82.480 116.590 82.740 ;
        RECT 116.650 82.480 116.910 82.740 ;
        RECT 116.970 82.480 117.230 82.740 ;
        RECT 117.290 82.480 117.550 82.740 ;
        RECT 117.610 82.480 117.870 82.740 ;
        RECT 138.525 82.480 138.785 82.740 ;
        RECT 138.845 82.480 139.105 82.740 ;
        RECT 139.165 82.480 139.425 82.740 ;
        RECT 139.485 82.480 139.745 82.740 ;
        RECT 139.805 82.480 140.065 82.740 ;
        RECT 60.845 79.760 61.105 80.020 ;
        RECT 61.165 79.760 61.425 80.020 ;
        RECT 61.485 79.760 61.745 80.020 ;
        RECT 61.805 79.760 62.065 80.020 ;
        RECT 62.125 79.760 62.385 80.020 ;
        RECT 83.040 79.760 83.300 80.020 ;
        RECT 83.360 79.760 83.620 80.020 ;
        RECT 83.680 79.760 83.940 80.020 ;
        RECT 84.000 79.760 84.260 80.020 ;
        RECT 84.320 79.760 84.580 80.020 ;
        RECT 105.235 79.760 105.495 80.020 ;
        RECT 105.555 79.760 105.815 80.020 ;
        RECT 105.875 79.760 106.135 80.020 ;
        RECT 106.195 79.760 106.455 80.020 ;
        RECT 106.515 79.760 106.775 80.020 ;
        RECT 127.430 79.760 127.690 80.020 ;
        RECT 127.750 79.760 128.010 80.020 ;
        RECT 128.070 79.760 128.330 80.020 ;
        RECT 128.390 79.760 128.650 80.020 ;
        RECT 128.710 79.760 128.970 80.020 ;
        RECT 71.940 77.040 72.200 77.300 ;
        RECT 72.260 77.040 72.520 77.300 ;
        RECT 72.580 77.040 72.840 77.300 ;
        RECT 72.900 77.040 73.160 77.300 ;
        RECT 73.220 77.040 73.480 77.300 ;
        RECT 94.135 77.040 94.395 77.300 ;
        RECT 94.455 77.040 94.715 77.300 ;
        RECT 94.775 77.040 95.035 77.300 ;
        RECT 95.095 77.040 95.355 77.300 ;
        RECT 95.415 77.040 95.675 77.300 ;
        RECT 116.330 77.040 116.590 77.300 ;
        RECT 116.650 77.040 116.910 77.300 ;
        RECT 116.970 77.040 117.230 77.300 ;
        RECT 117.290 77.040 117.550 77.300 ;
        RECT 117.610 77.040 117.870 77.300 ;
        RECT 138.525 77.040 138.785 77.300 ;
        RECT 138.845 77.040 139.105 77.300 ;
        RECT 139.165 77.040 139.425 77.300 ;
        RECT 139.485 77.040 139.745 77.300 ;
        RECT 139.805 77.040 140.065 77.300 ;
        RECT 60.845 74.320 61.105 74.580 ;
        RECT 61.165 74.320 61.425 74.580 ;
        RECT 61.485 74.320 61.745 74.580 ;
        RECT 61.805 74.320 62.065 74.580 ;
        RECT 62.125 74.320 62.385 74.580 ;
        RECT 83.040 74.320 83.300 74.580 ;
        RECT 83.360 74.320 83.620 74.580 ;
        RECT 83.680 74.320 83.940 74.580 ;
        RECT 84.000 74.320 84.260 74.580 ;
        RECT 84.320 74.320 84.580 74.580 ;
        RECT 105.235 74.320 105.495 74.580 ;
        RECT 105.555 74.320 105.815 74.580 ;
        RECT 105.875 74.320 106.135 74.580 ;
        RECT 106.195 74.320 106.455 74.580 ;
        RECT 106.515 74.320 106.775 74.580 ;
        RECT 127.430 74.320 127.690 74.580 ;
        RECT 127.750 74.320 128.010 74.580 ;
        RECT 128.070 74.320 128.330 74.580 ;
        RECT 128.390 74.320 128.650 74.580 ;
        RECT 128.710 74.320 128.970 74.580 ;
        RECT 71.940 71.600 72.200 71.860 ;
        RECT 72.260 71.600 72.520 71.860 ;
        RECT 72.580 71.600 72.840 71.860 ;
        RECT 72.900 71.600 73.160 71.860 ;
        RECT 73.220 71.600 73.480 71.860 ;
        RECT 94.135 71.600 94.395 71.860 ;
        RECT 94.455 71.600 94.715 71.860 ;
        RECT 94.775 71.600 95.035 71.860 ;
        RECT 95.095 71.600 95.355 71.860 ;
        RECT 95.415 71.600 95.675 71.860 ;
        RECT 116.330 71.600 116.590 71.860 ;
        RECT 116.650 71.600 116.910 71.860 ;
        RECT 116.970 71.600 117.230 71.860 ;
        RECT 117.290 71.600 117.550 71.860 ;
        RECT 117.610 71.600 117.870 71.860 ;
        RECT 138.525 71.600 138.785 71.860 ;
        RECT 138.845 71.600 139.105 71.860 ;
        RECT 139.165 71.600 139.425 71.860 ;
        RECT 139.485 71.600 139.745 71.860 ;
        RECT 139.805 71.600 140.065 71.860 ;
        RECT 60.845 68.880 61.105 69.140 ;
        RECT 61.165 68.880 61.425 69.140 ;
        RECT 61.485 68.880 61.745 69.140 ;
        RECT 61.805 68.880 62.065 69.140 ;
        RECT 62.125 68.880 62.385 69.140 ;
        RECT 83.040 68.880 83.300 69.140 ;
        RECT 83.360 68.880 83.620 69.140 ;
        RECT 83.680 68.880 83.940 69.140 ;
        RECT 84.000 68.880 84.260 69.140 ;
        RECT 84.320 68.880 84.580 69.140 ;
        RECT 105.235 68.880 105.495 69.140 ;
        RECT 105.555 68.880 105.815 69.140 ;
        RECT 105.875 68.880 106.135 69.140 ;
        RECT 106.195 68.880 106.455 69.140 ;
        RECT 106.515 68.880 106.775 69.140 ;
        RECT 127.430 68.880 127.690 69.140 ;
        RECT 127.750 68.880 128.010 69.140 ;
        RECT 128.070 68.880 128.330 69.140 ;
        RECT 128.390 68.880 128.650 69.140 ;
        RECT 128.710 68.880 128.970 69.140 ;
        RECT 71.940 66.160 72.200 66.420 ;
        RECT 72.260 66.160 72.520 66.420 ;
        RECT 72.580 66.160 72.840 66.420 ;
        RECT 72.900 66.160 73.160 66.420 ;
        RECT 73.220 66.160 73.480 66.420 ;
        RECT 94.135 66.160 94.395 66.420 ;
        RECT 94.455 66.160 94.715 66.420 ;
        RECT 94.775 66.160 95.035 66.420 ;
        RECT 95.095 66.160 95.355 66.420 ;
        RECT 95.415 66.160 95.675 66.420 ;
        RECT 116.330 66.160 116.590 66.420 ;
        RECT 116.650 66.160 116.910 66.420 ;
        RECT 116.970 66.160 117.230 66.420 ;
        RECT 117.290 66.160 117.550 66.420 ;
        RECT 117.610 66.160 117.870 66.420 ;
        RECT 138.525 66.160 138.785 66.420 ;
        RECT 138.845 66.160 139.105 66.420 ;
        RECT 139.165 66.160 139.425 66.420 ;
        RECT 139.485 66.160 139.745 66.420 ;
        RECT 139.805 66.160 140.065 66.420 ;
        RECT 60.845 63.440 61.105 63.700 ;
        RECT 61.165 63.440 61.425 63.700 ;
        RECT 61.485 63.440 61.745 63.700 ;
        RECT 61.805 63.440 62.065 63.700 ;
        RECT 62.125 63.440 62.385 63.700 ;
        RECT 83.040 63.440 83.300 63.700 ;
        RECT 83.360 63.440 83.620 63.700 ;
        RECT 83.680 63.440 83.940 63.700 ;
        RECT 84.000 63.440 84.260 63.700 ;
        RECT 84.320 63.440 84.580 63.700 ;
        RECT 105.235 63.440 105.495 63.700 ;
        RECT 105.555 63.440 105.815 63.700 ;
        RECT 105.875 63.440 106.135 63.700 ;
        RECT 106.195 63.440 106.455 63.700 ;
        RECT 106.515 63.440 106.775 63.700 ;
        RECT 127.430 63.440 127.690 63.700 ;
        RECT 127.750 63.440 128.010 63.700 ;
        RECT 128.070 63.440 128.330 63.700 ;
        RECT 128.390 63.440 128.650 63.700 ;
        RECT 128.710 63.440 128.970 63.700 ;
        RECT 71.940 60.720 72.200 60.980 ;
        RECT 72.260 60.720 72.520 60.980 ;
        RECT 72.580 60.720 72.840 60.980 ;
        RECT 72.900 60.720 73.160 60.980 ;
        RECT 73.220 60.720 73.480 60.980 ;
        RECT 94.135 60.720 94.395 60.980 ;
        RECT 94.455 60.720 94.715 60.980 ;
        RECT 94.775 60.720 95.035 60.980 ;
        RECT 95.095 60.720 95.355 60.980 ;
        RECT 95.415 60.720 95.675 60.980 ;
        RECT 116.330 60.720 116.590 60.980 ;
        RECT 116.650 60.720 116.910 60.980 ;
        RECT 116.970 60.720 117.230 60.980 ;
        RECT 117.290 60.720 117.550 60.980 ;
        RECT 117.610 60.720 117.870 60.980 ;
        RECT 138.525 60.720 138.785 60.980 ;
        RECT 138.845 60.720 139.105 60.980 ;
        RECT 139.165 60.720 139.425 60.980 ;
        RECT 139.485 60.720 139.745 60.980 ;
        RECT 139.805 60.720 140.065 60.980 ;
      LAYER met2 ;
        RECT 71.940 136.825 73.480 137.195 ;
        RECT 94.135 136.825 95.675 137.195 ;
        RECT 116.330 136.825 117.870 137.195 ;
        RECT 138.525 136.825 140.065 137.195 ;
        RECT 60.845 134.105 62.385 134.475 ;
        RECT 83.040 134.105 84.580 134.475 ;
        RECT 105.235 134.105 106.775 134.475 ;
        RECT 127.430 134.105 128.970 134.475 ;
        RECT 71.940 131.385 73.480 131.755 ;
        RECT 94.135 131.385 95.675 131.755 ;
        RECT 116.330 131.385 117.870 131.755 ;
        RECT 138.525 131.385 140.065 131.755 ;
        RECT 60.845 128.665 62.385 129.035 ;
        RECT 83.040 128.665 84.580 129.035 ;
        RECT 105.235 128.665 106.775 129.035 ;
        RECT 127.430 128.665 128.970 129.035 ;
        RECT 71.940 125.945 73.480 126.315 ;
        RECT 94.135 125.945 95.675 126.315 ;
        RECT 116.330 125.945 117.870 126.315 ;
        RECT 138.525 125.945 140.065 126.315 ;
        RECT 60.845 123.225 62.385 123.595 ;
        RECT 83.040 123.225 84.580 123.595 ;
        RECT 105.235 123.225 106.775 123.595 ;
        RECT 127.430 123.225 128.970 123.595 ;
        RECT 71.940 120.505 73.480 120.875 ;
        RECT 94.135 120.505 95.675 120.875 ;
        RECT 116.330 120.505 117.870 120.875 ;
        RECT 138.525 120.505 140.065 120.875 ;
        RECT 60.845 117.785 62.385 118.155 ;
        RECT 83.040 117.785 84.580 118.155 ;
        RECT 105.235 117.785 106.775 118.155 ;
        RECT 127.430 117.785 128.970 118.155 ;
        RECT 71.940 115.065 73.480 115.435 ;
        RECT 94.135 115.065 95.675 115.435 ;
        RECT 116.330 115.065 117.870 115.435 ;
        RECT 138.525 115.065 140.065 115.435 ;
        RECT 60.845 112.345 62.385 112.715 ;
        RECT 83.040 112.345 84.580 112.715 ;
        RECT 105.235 112.345 106.775 112.715 ;
        RECT 127.430 112.345 128.970 112.715 ;
        RECT 71.940 109.625 73.480 109.995 ;
        RECT 94.135 109.625 95.675 109.995 ;
        RECT 116.330 109.625 117.870 109.995 ;
        RECT 138.525 109.625 140.065 109.995 ;
        RECT 63.960 108.460 64.220 108.780 ;
        RECT 60.845 106.905 62.385 107.275 ;
        RECT 57.060 105.400 57.320 105.720 ;
        RECT 60.280 105.400 60.540 105.720 ;
        RECT 62.580 105.400 62.840 105.720 ;
        RECT 57.120 104.020 57.260 105.400 ;
        RECT 58.900 105.060 59.160 105.380 ;
        RECT 58.960 104.895 59.100 105.060 ;
        RECT 58.890 104.525 59.170 104.895 ;
        RECT 57.060 103.700 57.320 104.020 ;
        RECT 60.340 103.340 60.480 105.400 ;
        RECT 48.780 103.020 49.040 103.340 ;
        RECT 60.280 103.020 60.540 103.340 ;
        RECT 48.840 101.495 48.980 103.020 ;
        RECT 62.640 103.000 62.780 105.400 ;
        RECT 63.500 103.360 63.760 103.680 ;
        RECT 62.580 102.680 62.840 103.000 ;
        RECT 48.770 101.125 49.050 101.495 ;
        RECT 60.845 101.465 62.385 101.835 ;
        RECT 58.900 99.960 59.160 100.280 ;
        RECT 58.440 99.280 58.700 99.600 ;
        RECT 58.500 94.840 58.640 99.280 ;
        RECT 58.960 98.095 59.100 99.960 ;
        RECT 62.640 98.580 62.780 102.680 ;
        RECT 62.580 98.260 62.840 98.580 ;
        RECT 58.890 97.725 59.170 98.095 ;
        RECT 60.280 97.580 60.540 97.900 ;
        RECT 58.440 94.520 58.700 94.840 ;
        RECT 57.980 93.840 58.240 94.160 ;
        RECT 58.040 93.140 58.180 93.840 ;
        RECT 58.500 93.140 58.640 94.520 ;
        RECT 60.340 93.140 60.480 97.580 ;
        RECT 60.845 96.025 62.385 96.395 ;
        RECT 57.980 92.820 58.240 93.140 ;
        RECT 58.440 92.820 58.700 93.140 ;
        RECT 60.280 92.820 60.540 93.140 ;
        RECT 58.500 91.860 58.640 92.820 ;
        RECT 62.580 92.140 62.840 92.460 ;
        RECT 58.500 91.720 59.100 91.860 ;
        RECT 58.960 89.740 59.100 91.720 ;
        RECT 60.280 91.120 60.540 91.440 ;
        RECT 58.900 89.420 59.160 89.740 ;
        RECT 60.340 89.400 60.480 91.120 ;
        RECT 60.845 90.585 62.385 90.955 ;
        RECT 62.640 90.420 62.780 92.140 ;
        RECT 63.560 92.120 63.700 103.360 ;
        RECT 64.020 103.000 64.160 108.460 ;
        RECT 83.040 106.905 84.580 107.275 ;
        RECT 105.235 106.905 106.775 107.275 ;
        RECT 127.430 106.905 128.970 107.275 ;
        RECT 71.940 104.185 73.480 104.555 ;
        RECT 94.135 104.185 95.675 104.555 ;
        RECT 116.330 104.185 117.870 104.555 ;
        RECT 138.525 104.185 140.065 104.555 ;
        RECT 63.960 102.680 64.220 103.000 ;
        RECT 64.020 94.840 64.160 102.680 ;
        RECT 83.040 101.465 84.580 101.835 ;
        RECT 105.235 101.465 106.775 101.835 ;
        RECT 127.430 101.465 128.970 101.835 ;
        RECT 71.940 98.745 73.480 99.115 ;
        RECT 94.135 98.745 95.675 99.115 ;
        RECT 116.330 98.745 117.870 99.115 ;
        RECT 138.525 98.745 140.065 99.115 ;
        RECT 83.040 96.025 84.580 96.395 ;
        RECT 105.235 96.025 106.775 96.395 ;
        RECT 127.430 96.025 128.970 96.395 ;
        RECT 63.960 94.520 64.220 94.840 ;
        RECT 66.260 93.840 66.520 94.160 ;
        RECT 66.320 92.460 66.460 93.840 ;
        RECT 71.940 93.305 73.480 93.675 ;
        RECT 94.135 93.305 95.675 93.675 ;
        RECT 116.330 93.305 117.870 93.675 ;
        RECT 138.525 93.305 140.065 93.675 ;
        RECT 66.260 92.140 66.520 92.460 ;
        RECT 63.500 91.800 63.760 92.120 ;
        RECT 83.040 90.585 84.580 90.955 ;
        RECT 105.235 90.585 106.775 90.955 ;
        RECT 127.430 90.585 128.970 90.955 ;
        RECT 62.580 90.100 62.840 90.420 ;
        RECT 60.280 89.080 60.540 89.400 ;
        RECT 71.940 87.865 73.480 88.235 ;
        RECT 94.135 87.865 95.675 88.235 ;
        RECT 116.330 87.865 117.870 88.235 ;
        RECT 138.525 87.865 140.065 88.235 ;
        RECT 60.845 85.145 62.385 85.515 ;
        RECT 83.040 85.145 84.580 85.515 ;
        RECT 105.235 85.145 106.775 85.515 ;
        RECT 127.430 85.145 128.970 85.515 ;
        RECT 71.940 82.425 73.480 82.795 ;
        RECT 94.135 82.425 95.675 82.795 ;
        RECT 116.330 82.425 117.870 82.795 ;
        RECT 138.525 82.425 140.065 82.795 ;
        RECT 60.845 79.705 62.385 80.075 ;
        RECT 83.040 79.705 84.580 80.075 ;
        RECT 105.235 79.705 106.775 80.075 ;
        RECT 127.430 79.705 128.970 80.075 ;
        RECT 71.940 76.985 73.480 77.355 ;
        RECT 94.135 76.985 95.675 77.355 ;
        RECT 116.330 76.985 117.870 77.355 ;
        RECT 138.525 76.985 140.065 77.355 ;
        RECT 60.845 74.265 62.385 74.635 ;
        RECT 83.040 74.265 84.580 74.635 ;
        RECT 105.235 74.265 106.775 74.635 ;
        RECT 127.430 74.265 128.970 74.635 ;
        RECT 71.940 71.545 73.480 71.915 ;
        RECT 94.135 71.545 95.675 71.915 ;
        RECT 116.330 71.545 117.870 71.915 ;
        RECT 138.525 71.545 140.065 71.915 ;
        RECT 60.845 68.825 62.385 69.195 ;
        RECT 83.040 68.825 84.580 69.195 ;
        RECT 105.235 68.825 106.775 69.195 ;
        RECT 127.430 68.825 128.970 69.195 ;
        RECT 71.940 66.105 73.480 66.475 ;
        RECT 94.135 66.105 95.675 66.475 ;
        RECT 116.330 66.105 117.870 66.475 ;
        RECT 138.525 66.105 140.065 66.475 ;
        RECT 60.845 63.385 62.385 63.755 ;
        RECT 83.040 63.385 84.580 63.755 ;
        RECT 105.235 63.385 106.775 63.755 ;
        RECT 127.430 63.385 128.970 63.755 ;
        RECT 71.940 60.665 73.480 61.035 ;
        RECT 94.135 60.665 95.675 61.035 ;
        RECT 116.330 60.665 117.870 61.035 ;
        RECT 138.525 60.665 140.065 61.035 ;
      LAYER via2 ;
        RECT 71.970 136.870 72.250 137.150 ;
        RECT 72.370 136.870 72.650 137.150 ;
        RECT 72.770 136.870 73.050 137.150 ;
        RECT 73.170 136.870 73.450 137.150 ;
        RECT 94.165 136.870 94.445 137.150 ;
        RECT 94.565 136.870 94.845 137.150 ;
        RECT 94.965 136.870 95.245 137.150 ;
        RECT 95.365 136.870 95.645 137.150 ;
        RECT 116.360 136.870 116.640 137.150 ;
        RECT 116.760 136.870 117.040 137.150 ;
        RECT 117.160 136.870 117.440 137.150 ;
        RECT 117.560 136.870 117.840 137.150 ;
        RECT 138.555 136.870 138.835 137.150 ;
        RECT 138.955 136.870 139.235 137.150 ;
        RECT 139.355 136.870 139.635 137.150 ;
        RECT 139.755 136.870 140.035 137.150 ;
        RECT 60.875 134.150 61.155 134.430 ;
        RECT 61.275 134.150 61.555 134.430 ;
        RECT 61.675 134.150 61.955 134.430 ;
        RECT 62.075 134.150 62.355 134.430 ;
        RECT 83.070 134.150 83.350 134.430 ;
        RECT 83.470 134.150 83.750 134.430 ;
        RECT 83.870 134.150 84.150 134.430 ;
        RECT 84.270 134.150 84.550 134.430 ;
        RECT 105.265 134.150 105.545 134.430 ;
        RECT 105.665 134.150 105.945 134.430 ;
        RECT 106.065 134.150 106.345 134.430 ;
        RECT 106.465 134.150 106.745 134.430 ;
        RECT 127.460 134.150 127.740 134.430 ;
        RECT 127.860 134.150 128.140 134.430 ;
        RECT 128.260 134.150 128.540 134.430 ;
        RECT 128.660 134.150 128.940 134.430 ;
        RECT 71.970 131.430 72.250 131.710 ;
        RECT 72.370 131.430 72.650 131.710 ;
        RECT 72.770 131.430 73.050 131.710 ;
        RECT 73.170 131.430 73.450 131.710 ;
        RECT 94.165 131.430 94.445 131.710 ;
        RECT 94.565 131.430 94.845 131.710 ;
        RECT 94.965 131.430 95.245 131.710 ;
        RECT 95.365 131.430 95.645 131.710 ;
        RECT 116.360 131.430 116.640 131.710 ;
        RECT 116.760 131.430 117.040 131.710 ;
        RECT 117.160 131.430 117.440 131.710 ;
        RECT 117.560 131.430 117.840 131.710 ;
        RECT 138.555 131.430 138.835 131.710 ;
        RECT 138.955 131.430 139.235 131.710 ;
        RECT 139.355 131.430 139.635 131.710 ;
        RECT 139.755 131.430 140.035 131.710 ;
        RECT 60.875 128.710 61.155 128.990 ;
        RECT 61.275 128.710 61.555 128.990 ;
        RECT 61.675 128.710 61.955 128.990 ;
        RECT 62.075 128.710 62.355 128.990 ;
        RECT 83.070 128.710 83.350 128.990 ;
        RECT 83.470 128.710 83.750 128.990 ;
        RECT 83.870 128.710 84.150 128.990 ;
        RECT 84.270 128.710 84.550 128.990 ;
        RECT 105.265 128.710 105.545 128.990 ;
        RECT 105.665 128.710 105.945 128.990 ;
        RECT 106.065 128.710 106.345 128.990 ;
        RECT 106.465 128.710 106.745 128.990 ;
        RECT 127.460 128.710 127.740 128.990 ;
        RECT 127.860 128.710 128.140 128.990 ;
        RECT 128.260 128.710 128.540 128.990 ;
        RECT 128.660 128.710 128.940 128.990 ;
        RECT 71.970 125.990 72.250 126.270 ;
        RECT 72.370 125.990 72.650 126.270 ;
        RECT 72.770 125.990 73.050 126.270 ;
        RECT 73.170 125.990 73.450 126.270 ;
        RECT 94.165 125.990 94.445 126.270 ;
        RECT 94.565 125.990 94.845 126.270 ;
        RECT 94.965 125.990 95.245 126.270 ;
        RECT 95.365 125.990 95.645 126.270 ;
        RECT 116.360 125.990 116.640 126.270 ;
        RECT 116.760 125.990 117.040 126.270 ;
        RECT 117.160 125.990 117.440 126.270 ;
        RECT 117.560 125.990 117.840 126.270 ;
        RECT 138.555 125.990 138.835 126.270 ;
        RECT 138.955 125.990 139.235 126.270 ;
        RECT 139.355 125.990 139.635 126.270 ;
        RECT 139.755 125.990 140.035 126.270 ;
        RECT 60.875 123.270 61.155 123.550 ;
        RECT 61.275 123.270 61.555 123.550 ;
        RECT 61.675 123.270 61.955 123.550 ;
        RECT 62.075 123.270 62.355 123.550 ;
        RECT 83.070 123.270 83.350 123.550 ;
        RECT 83.470 123.270 83.750 123.550 ;
        RECT 83.870 123.270 84.150 123.550 ;
        RECT 84.270 123.270 84.550 123.550 ;
        RECT 105.265 123.270 105.545 123.550 ;
        RECT 105.665 123.270 105.945 123.550 ;
        RECT 106.065 123.270 106.345 123.550 ;
        RECT 106.465 123.270 106.745 123.550 ;
        RECT 127.460 123.270 127.740 123.550 ;
        RECT 127.860 123.270 128.140 123.550 ;
        RECT 128.260 123.270 128.540 123.550 ;
        RECT 128.660 123.270 128.940 123.550 ;
        RECT 71.970 120.550 72.250 120.830 ;
        RECT 72.370 120.550 72.650 120.830 ;
        RECT 72.770 120.550 73.050 120.830 ;
        RECT 73.170 120.550 73.450 120.830 ;
        RECT 94.165 120.550 94.445 120.830 ;
        RECT 94.565 120.550 94.845 120.830 ;
        RECT 94.965 120.550 95.245 120.830 ;
        RECT 95.365 120.550 95.645 120.830 ;
        RECT 116.360 120.550 116.640 120.830 ;
        RECT 116.760 120.550 117.040 120.830 ;
        RECT 117.160 120.550 117.440 120.830 ;
        RECT 117.560 120.550 117.840 120.830 ;
        RECT 138.555 120.550 138.835 120.830 ;
        RECT 138.955 120.550 139.235 120.830 ;
        RECT 139.355 120.550 139.635 120.830 ;
        RECT 139.755 120.550 140.035 120.830 ;
        RECT 60.875 117.830 61.155 118.110 ;
        RECT 61.275 117.830 61.555 118.110 ;
        RECT 61.675 117.830 61.955 118.110 ;
        RECT 62.075 117.830 62.355 118.110 ;
        RECT 83.070 117.830 83.350 118.110 ;
        RECT 83.470 117.830 83.750 118.110 ;
        RECT 83.870 117.830 84.150 118.110 ;
        RECT 84.270 117.830 84.550 118.110 ;
        RECT 105.265 117.830 105.545 118.110 ;
        RECT 105.665 117.830 105.945 118.110 ;
        RECT 106.065 117.830 106.345 118.110 ;
        RECT 106.465 117.830 106.745 118.110 ;
        RECT 127.460 117.830 127.740 118.110 ;
        RECT 127.860 117.830 128.140 118.110 ;
        RECT 128.260 117.830 128.540 118.110 ;
        RECT 128.660 117.830 128.940 118.110 ;
        RECT 71.970 115.110 72.250 115.390 ;
        RECT 72.370 115.110 72.650 115.390 ;
        RECT 72.770 115.110 73.050 115.390 ;
        RECT 73.170 115.110 73.450 115.390 ;
        RECT 94.165 115.110 94.445 115.390 ;
        RECT 94.565 115.110 94.845 115.390 ;
        RECT 94.965 115.110 95.245 115.390 ;
        RECT 95.365 115.110 95.645 115.390 ;
        RECT 116.360 115.110 116.640 115.390 ;
        RECT 116.760 115.110 117.040 115.390 ;
        RECT 117.160 115.110 117.440 115.390 ;
        RECT 117.560 115.110 117.840 115.390 ;
        RECT 138.555 115.110 138.835 115.390 ;
        RECT 138.955 115.110 139.235 115.390 ;
        RECT 139.355 115.110 139.635 115.390 ;
        RECT 139.755 115.110 140.035 115.390 ;
        RECT 60.875 112.390 61.155 112.670 ;
        RECT 61.275 112.390 61.555 112.670 ;
        RECT 61.675 112.390 61.955 112.670 ;
        RECT 62.075 112.390 62.355 112.670 ;
        RECT 83.070 112.390 83.350 112.670 ;
        RECT 83.470 112.390 83.750 112.670 ;
        RECT 83.870 112.390 84.150 112.670 ;
        RECT 84.270 112.390 84.550 112.670 ;
        RECT 105.265 112.390 105.545 112.670 ;
        RECT 105.665 112.390 105.945 112.670 ;
        RECT 106.065 112.390 106.345 112.670 ;
        RECT 106.465 112.390 106.745 112.670 ;
        RECT 127.460 112.390 127.740 112.670 ;
        RECT 127.860 112.390 128.140 112.670 ;
        RECT 128.260 112.390 128.540 112.670 ;
        RECT 128.660 112.390 128.940 112.670 ;
        RECT 71.970 109.670 72.250 109.950 ;
        RECT 72.370 109.670 72.650 109.950 ;
        RECT 72.770 109.670 73.050 109.950 ;
        RECT 73.170 109.670 73.450 109.950 ;
        RECT 94.165 109.670 94.445 109.950 ;
        RECT 94.565 109.670 94.845 109.950 ;
        RECT 94.965 109.670 95.245 109.950 ;
        RECT 95.365 109.670 95.645 109.950 ;
        RECT 116.360 109.670 116.640 109.950 ;
        RECT 116.760 109.670 117.040 109.950 ;
        RECT 117.160 109.670 117.440 109.950 ;
        RECT 117.560 109.670 117.840 109.950 ;
        RECT 138.555 109.670 138.835 109.950 ;
        RECT 138.955 109.670 139.235 109.950 ;
        RECT 139.355 109.670 139.635 109.950 ;
        RECT 139.755 109.670 140.035 109.950 ;
        RECT 60.875 106.950 61.155 107.230 ;
        RECT 61.275 106.950 61.555 107.230 ;
        RECT 61.675 106.950 61.955 107.230 ;
        RECT 62.075 106.950 62.355 107.230 ;
        RECT 58.890 104.570 59.170 104.850 ;
        RECT 60.875 101.510 61.155 101.790 ;
        RECT 61.275 101.510 61.555 101.790 ;
        RECT 61.675 101.510 61.955 101.790 ;
        RECT 62.075 101.510 62.355 101.790 ;
        RECT 48.770 101.170 49.050 101.450 ;
        RECT 58.890 97.770 59.170 98.050 ;
        RECT 60.875 96.070 61.155 96.350 ;
        RECT 61.275 96.070 61.555 96.350 ;
        RECT 61.675 96.070 61.955 96.350 ;
        RECT 62.075 96.070 62.355 96.350 ;
        RECT 60.875 90.630 61.155 90.910 ;
        RECT 61.275 90.630 61.555 90.910 ;
        RECT 61.675 90.630 61.955 90.910 ;
        RECT 62.075 90.630 62.355 90.910 ;
        RECT 83.070 106.950 83.350 107.230 ;
        RECT 83.470 106.950 83.750 107.230 ;
        RECT 83.870 106.950 84.150 107.230 ;
        RECT 84.270 106.950 84.550 107.230 ;
        RECT 105.265 106.950 105.545 107.230 ;
        RECT 105.665 106.950 105.945 107.230 ;
        RECT 106.065 106.950 106.345 107.230 ;
        RECT 106.465 106.950 106.745 107.230 ;
        RECT 127.460 106.950 127.740 107.230 ;
        RECT 127.860 106.950 128.140 107.230 ;
        RECT 128.260 106.950 128.540 107.230 ;
        RECT 128.660 106.950 128.940 107.230 ;
        RECT 71.970 104.230 72.250 104.510 ;
        RECT 72.370 104.230 72.650 104.510 ;
        RECT 72.770 104.230 73.050 104.510 ;
        RECT 73.170 104.230 73.450 104.510 ;
        RECT 94.165 104.230 94.445 104.510 ;
        RECT 94.565 104.230 94.845 104.510 ;
        RECT 94.965 104.230 95.245 104.510 ;
        RECT 95.365 104.230 95.645 104.510 ;
        RECT 116.360 104.230 116.640 104.510 ;
        RECT 116.760 104.230 117.040 104.510 ;
        RECT 117.160 104.230 117.440 104.510 ;
        RECT 117.560 104.230 117.840 104.510 ;
        RECT 138.555 104.230 138.835 104.510 ;
        RECT 138.955 104.230 139.235 104.510 ;
        RECT 139.355 104.230 139.635 104.510 ;
        RECT 139.755 104.230 140.035 104.510 ;
        RECT 83.070 101.510 83.350 101.790 ;
        RECT 83.470 101.510 83.750 101.790 ;
        RECT 83.870 101.510 84.150 101.790 ;
        RECT 84.270 101.510 84.550 101.790 ;
        RECT 105.265 101.510 105.545 101.790 ;
        RECT 105.665 101.510 105.945 101.790 ;
        RECT 106.065 101.510 106.345 101.790 ;
        RECT 106.465 101.510 106.745 101.790 ;
        RECT 127.460 101.510 127.740 101.790 ;
        RECT 127.860 101.510 128.140 101.790 ;
        RECT 128.260 101.510 128.540 101.790 ;
        RECT 128.660 101.510 128.940 101.790 ;
        RECT 71.970 98.790 72.250 99.070 ;
        RECT 72.370 98.790 72.650 99.070 ;
        RECT 72.770 98.790 73.050 99.070 ;
        RECT 73.170 98.790 73.450 99.070 ;
        RECT 94.165 98.790 94.445 99.070 ;
        RECT 94.565 98.790 94.845 99.070 ;
        RECT 94.965 98.790 95.245 99.070 ;
        RECT 95.365 98.790 95.645 99.070 ;
        RECT 116.360 98.790 116.640 99.070 ;
        RECT 116.760 98.790 117.040 99.070 ;
        RECT 117.160 98.790 117.440 99.070 ;
        RECT 117.560 98.790 117.840 99.070 ;
        RECT 138.555 98.790 138.835 99.070 ;
        RECT 138.955 98.790 139.235 99.070 ;
        RECT 139.355 98.790 139.635 99.070 ;
        RECT 139.755 98.790 140.035 99.070 ;
        RECT 83.070 96.070 83.350 96.350 ;
        RECT 83.470 96.070 83.750 96.350 ;
        RECT 83.870 96.070 84.150 96.350 ;
        RECT 84.270 96.070 84.550 96.350 ;
        RECT 105.265 96.070 105.545 96.350 ;
        RECT 105.665 96.070 105.945 96.350 ;
        RECT 106.065 96.070 106.345 96.350 ;
        RECT 106.465 96.070 106.745 96.350 ;
        RECT 127.460 96.070 127.740 96.350 ;
        RECT 127.860 96.070 128.140 96.350 ;
        RECT 128.260 96.070 128.540 96.350 ;
        RECT 128.660 96.070 128.940 96.350 ;
        RECT 71.970 93.350 72.250 93.630 ;
        RECT 72.370 93.350 72.650 93.630 ;
        RECT 72.770 93.350 73.050 93.630 ;
        RECT 73.170 93.350 73.450 93.630 ;
        RECT 94.165 93.350 94.445 93.630 ;
        RECT 94.565 93.350 94.845 93.630 ;
        RECT 94.965 93.350 95.245 93.630 ;
        RECT 95.365 93.350 95.645 93.630 ;
        RECT 116.360 93.350 116.640 93.630 ;
        RECT 116.760 93.350 117.040 93.630 ;
        RECT 117.160 93.350 117.440 93.630 ;
        RECT 117.560 93.350 117.840 93.630 ;
        RECT 138.555 93.350 138.835 93.630 ;
        RECT 138.955 93.350 139.235 93.630 ;
        RECT 139.355 93.350 139.635 93.630 ;
        RECT 139.755 93.350 140.035 93.630 ;
        RECT 83.070 90.630 83.350 90.910 ;
        RECT 83.470 90.630 83.750 90.910 ;
        RECT 83.870 90.630 84.150 90.910 ;
        RECT 84.270 90.630 84.550 90.910 ;
        RECT 105.265 90.630 105.545 90.910 ;
        RECT 105.665 90.630 105.945 90.910 ;
        RECT 106.065 90.630 106.345 90.910 ;
        RECT 106.465 90.630 106.745 90.910 ;
        RECT 127.460 90.630 127.740 90.910 ;
        RECT 127.860 90.630 128.140 90.910 ;
        RECT 128.260 90.630 128.540 90.910 ;
        RECT 128.660 90.630 128.940 90.910 ;
        RECT 71.970 87.910 72.250 88.190 ;
        RECT 72.370 87.910 72.650 88.190 ;
        RECT 72.770 87.910 73.050 88.190 ;
        RECT 73.170 87.910 73.450 88.190 ;
        RECT 94.165 87.910 94.445 88.190 ;
        RECT 94.565 87.910 94.845 88.190 ;
        RECT 94.965 87.910 95.245 88.190 ;
        RECT 95.365 87.910 95.645 88.190 ;
        RECT 116.360 87.910 116.640 88.190 ;
        RECT 116.760 87.910 117.040 88.190 ;
        RECT 117.160 87.910 117.440 88.190 ;
        RECT 117.560 87.910 117.840 88.190 ;
        RECT 138.555 87.910 138.835 88.190 ;
        RECT 138.955 87.910 139.235 88.190 ;
        RECT 139.355 87.910 139.635 88.190 ;
        RECT 139.755 87.910 140.035 88.190 ;
        RECT 60.875 85.190 61.155 85.470 ;
        RECT 61.275 85.190 61.555 85.470 ;
        RECT 61.675 85.190 61.955 85.470 ;
        RECT 62.075 85.190 62.355 85.470 ;
        RECT 83.070 85.190 83.350 85.470 ;
        RECT 83.470 85.190 83.750 85.470 ;
        RECT 83.870 85.190 84.150 85.470 ;
        RECT 84.270 85.190 84.550 85.470 ;
        RECT 105.265 85.190 105.545 85.470 ;
        RECT 105.665 85.190 105.945 85.470 ;
        RECT 106.065 85.190 106.345 85.470 ;
        RECT 106.465 85.190 106.745 85.470 ;
        RECT 127.460 85.190 127.740 85.470 ;
        RECT 127.860 85.190 128.140 85.470 ;
        RECT 128.260 85.190 128.540 85.470 ;
        RECT 128.660 85.190 128.940 85.470 ;
        RECT 71.970 82.470 72.250 82.750 ;
        RECT 72.370 82.470 72.650 82.750 ;
        RECT 72.770 82.470 73.050 82.750 ;
        RECT 73.170 82.470 73.450 82.750 ;
        RECT 94.165 82.470 94.445 82.750 ;
        RECT 94.565 82.470 94.845 82.750 ;
        RECT 94.965 82.470 95.245 82.750 ;
        RECT 95.365 82.470 95.645 82.750 ;
        RECT 116.360 82.470 116.640 82.750 ;
        RECT 116.760 82.470 117.040 82.750 ;
        RECT 117.160 82.470 117.440 82.750 ;
        RECT 117.560 82.470 117.840 82.750 ;
        RECT 138.555 82.470 138.835 82.750 ;
        RECT 138.955 82.470 139.235 82.750 ;
        RECT 139.355 82.470 139.635 82.750 ;
        RECT 139.755 82.470 140.035 82.750 ;
        RECT 60.875 79.750 61.155 80.030 ;
        RECT 61.275 79.750 61.555 80.030 ;
        RECT 61.675 79.750 61.955 80.030 ;
        RECT 62.075 79.750 62.355 80.030 ;
        RECT 83.070 79.750 83.350 80.030 ;
        RECT 83.470 79.750 83.750 80.030 ;
        RECT 83.870 79.750 84.150 80.030 ;
        RECT 84.270 79.750 84.550 80.030 ;
        RECT 105.265 79.750 105.545 80.030 ;
        RECT 105.665 79.750 105.945 80.030 ;
        RECT 106.065 79.750 106.345 80.030 ;
        RECT 106.465 79.750 106.745 80.030 ;
        RECT 127.460 79.750 127.740 80.030 ;
        RECT 127.860 79.750 128.140 80.030 ;
        RECT 128.260 79.750 128.540 80.030 ;
        RECT 128.660 79.750 128.940 80.030 ;
        RECT 71.970 77.030 72.250 77.310 ;
        RECT 72.370 77.030 72.650 77.310 ;
        RECT 72.770 77.030 73.050 77.310 ;
        RECT 73.170 77.030 73.450 77.310 ;
        RECT 94.165 77.030 94.445 77.310 ;
        RECT 94.565 77.030 94.845 77.310 ;
        RECT 94.965 77.030 95.245 77.310 ;
        RECT 95.365 77.030 95.645 77.310 ;
        RECT 116.360 77.030 116.640 77.310 ;
        RECT 116.760 77.030 117.040 77.310 ;
        RECT 117.160 77.030 117.440 77.310 ;
        RECT 117.560 77.030 117.840 77.310 ;
        RECT 138.555 77.030 138.835 77.310 ;
        RECT 138.955 77.030 139.235 77.310 ;
        RECT 139.355 77.030 139.635 77.310 ;
        RECT 139.755 77.030 140.035 77.310 ;
        RECT 60.875 74.310 61.155 74.590 ;
        RECT 61.275 74.310 61.555 74.590 ;
        RECT 61.675 74.310 61.955 74.590 ;
        RECT 62.075 74.310 62.355 74.590 ;
        RECT 83.070 74.310 83.350 74.590 ;
        RECT 83.470 74.310 83.750 74.590 ;
        RECT 83.870 74.310 84.150 74.590 ;
        RECT 84.270 74.310 84.550 74.590 ;
        RECT 105.265 74.310 105.545 74.590 ;
        RECT 105.665 74.310 105.945 74.590 ;
        RECT 106.065 74.310 106.345 74.590 ;
        RECT 106.465 74.310 106.745 74.590 ;
        RECT 127.460 74.310 127.740 74.590 ;
        RECT 127.860 74.310 128.140 74.590 ;
        RECT 128.260 74.310 128.540 74.590 ;
        RECT 128.660 74.310 128.940 74.590 ;
        RECT 71.970 71.590 72.250 71.870 ;
        RECT 72.370 71.590 72.650 71.870 ;
        RECT 72.770 71.590 73.050 71.870 ;
        RECT 73.170 71.590 73.450 71.870 ;
        RECT 94.165 71.590 94.445 71.870 ;
        RECT 94.565 71.590 94.845 71.870 ;
        RECT 94.965 71.590 95.245 71.870 ;
        RECT 95.365 71.590 95.645 71.870 ;
        RECT 116.360 71.590 116.640 71.870 ;
        RECT 116.760 71.590 117.040 71.870 ;
        RECT 117.160 71.590 117.440 71.870 ;
        RECT 117.560 71.590 117.840 71.870 ;
        RECT 138.555 71.590 138.835 71.870 ;
        RECT 138.955 71.590 139.235 71.870 ;
        RECT 139.355 71.590 139.635 71.870 ;
        RECT 139.755 71.590 140.035 71.870 ;
        RECT 60.875 68.870 61.155 69.150 ;
        RECT 61.275 68.870 61.555 69.150 ;
        RECT 61.675 68.870 61.955 69.150 ;
        RECT 62.075 68.870 62.355 69.150 ;
        RECT 83.070 68.870 83.350 69.150 ;
        RECT 83.470 68.870 83.750 69.150 ;
        RECT 83.870 68.870 84.150 69.150 ;
        RECT 84.270 68.870 84.550 69.150 ;
        RECT 105.265 68.870 105.545 69.150 ;
        RECT 105.665 68.870 105.945 69.150 ;
        RECT 106.065 68.870 106.345 69.150 ;
        RECT 106.465 68.870 106.745 69.150 ;
        RECT 127.460 68.870 127.740 69.150 ;
        RECT 127.860 68.870 128.140 69.150 ;
        RECT 128.260 68.870 128.540 69.150 ;
        RECT 128.660 68.870 128.940 69.150 ;
        RECT 71.970 66.150 72.250 66.430 ;
        RECT 72.370 66.150 72.650 66.430 ;
        RECT 72.770 66.150 73.050 66.430 ;
        RECT 73.170 66.150 73.450 66.430 ;
        RECT 94.165 66.150 94.445 66.430 ;
        RECT 94.565 66.150 94.845 66.430 ;
        RECT 94.965 66.150 95.245 66.430 ;
        RECT 95.365 66.150 95.645 66.430 ;
        RECT 116.360 66.150 116.640 66.430 ;
        RECT 116.760 66.150 117.040 66.430 ;
        RECT 117.160 66.150 117.440 66.430 ;
        RECT 117.560 66.150 117.840 66.430 ;
        RECT 138.555 66.150 138.835 66.430 ;
        RECT 138.955 66.150 139.235 66.430 ;
        RECT 139.355 66.150 139.635 66.430 ;
        RECT 139.755 66.150 140.035 66.430 ;
        RECT 60.875 63.430 61.155 63.710 ;
        RECT 61.275 63.430 61.555 63.710 ;
        RECT 61.675 63.430 61.955 63.710 ;
        RECT 62.075 63.430 62.355 63.710 ;
        RECT 83.070 63.430 83.350 63.710 ;
        RECT 83.470 63.430 83.750 63.710 ;
        RECT 83.870 63.430 84.150 63.710 ;
        RECT 84.270 63.430 84.550 63.710 ;
        RECT 105.265 63.430 105.545 63.710 ;
        RECT 105.665 63.430 105.945 63.710 ;
        RECT 106.065 63.430 106.345 63.710 ;
        RECT 106.465 63.430 106.745 63.710 ;
        RECT 127.460 63.430 127.740 63.710 ;
        RECT 127.860 63.430 128.140 63.710 ;
        RECT 128.260 63.430 128.540 63.710 ;
        RECT 128.660 63.430 128.940 63.710 ;
        RECT 71.970 60.710 72.250 60.990 ;
        RECT 72.370 60.710 72.650 60.990 ;
        RECT 72.770 60.710 73.050 60.990 ;
        RECT 73.170 60.710 73.450 60.990 ;
        RECT 94.165 60.710 94.445 60.990 ;
        RECT 94.565 60.710 94.845 60.990 ;
        RECT 94.965 60.710 95.245 60.990 ;
        RECT 95.365 60.710 95.645 60.990 ;
        RECT 116.360 60.710 116.640 60.990 ;
        RECT 116.760 60.710 117.040 60.990 ;
        RECT 117.160 60.710 117.440 60.990 ;
        RECT 117.560 60.710 117.840 60.990 ;
        RECT 138.555 60.710 138.835 60.990 ;
        RECT 138.955 60.710 139.235 60.990 ;
        RECT 139.355 60.710 139.635 60.990 ;
        RECT 139.755 60.710 140.035 60.990 ;
      LAYER met3 ;
        RECT 71.920 136.845 73.500 137.175 ;
        RECT 94.115 136.845 95.695 137.175 ;
        RECT 116.310 136.845 117.890 137.175 ;
        RECT 138.505 136.845 140.085 137.175 ;
        RECT 60.825 134.125 62.405 134.455 ;
        RECT 83.020 134.125 84.600 134.455 ;
        RECT 105.215 134.125 106.795 134.455 ;
        RECT 127.410 134.125 128.990 134.455 ;
        RECT 71.920 131.405 73.500 131.735 ;
        RECT 94.115 131.405 95.695 131.735 ;
        RECT 116.310 131.405 117.890 131.735 ;
        RECT 138.505 131.405 140.085 131.735 ;
        RECT 60.825 128.685 62.405 129.015 ;
        RECT 83.020 128.685 84.600 129.015 ;
        RECT 105.215 128.685 106.795 129.015 ;
        RECT 127.410 128.685 128.990 129.015 ;
        RECT 71.920 125.965 73.500 126.295 ;
        RECT 94.115 125.965 95.695 126.295 ;
        RECT 116.310 125.965 117.890 126.295 ;
        RECT 138.505 125.965 140.085 126.295 ;
        RECT 60.825 123.245 62.405 123.575 ;
        RECT 83.020 123.245 84.600 123.575 ;
        RECT 105.215 123.245 106.795 123.575 ;
        RECT 127.410 123.245 128.990 123.575 ;
        RECT 71.920 120.525 73.500 120.855 ;
        RECT 94.115 120.525 95.695 120.855 ;
        RECT 116.310 120.525 117.890 120.855 ;
        RECT 138.505 120.525 140.085 120.855 ;
        RECT 60.825 117.805 62.405 118.135 ;
        RECT 83.020 117.805 84.600 118.135 ;
        RECT 105.215 117.805 106.795 118.135 ;
        RECT 127.410 117.805 128.990 118.135 ;
        RECT 71.920 115.085 73.500 115.415 ;
        RECT 94.115 115.085 95.695 115.415 ;
        RECT 116.310 115.085 117.890 115.415 ;
        RECT 138.505 115.085 140.085 115.415 ;
        RECT 60.825 112.365 62.405 112.695 ;
        RECT 83.020 112.365 84.600 112.695 ;
        RECT 105.215 112.365 106.795 112.695 ;
        RECT 127.410 112.365 128.990 112.695 ;
        RECT 71.920 109.645 73.500 109.975 ;
        RECT 94.115 109.645 95.695 109.975 ;
        RECT 116.310 109.645 117.890 109.975 ;
        RECT 138.505 109.645 140.085 109.975 ;
        RECT 60.825 106.925 62.405 107.255 ;
        RECT 83.020 106.925 84.600 107.255 ;
        RECT 105.215 106.925 106.795 107.255 ;
        RECT 127.410 106.925 128.990 107.255 ;
        RECT 37.160 105.110 38.060 105.160 ;
        RECT 37.160 105.010 38.720 105.110 ;
        RECT 35.230 104.860 47.000 105.010 ;
        RECT 58.865 104.860 59.195 104.875 ;
        RECT 35.230 104.560 59.195 104.860 ;
        RECT 35.230 104.410 47.000 104.560 ;
        RECT 58.865 104.545 59.195 104.560 ;
        RECT 37.160 104.260 38.720 104.410 ;
        RECT 37.820 104.210 38.720 104.260 ;
        RECT 71.920 104.205 73.500 104.535 ;
        RECT 94.115 104.205 95.695 104.535 ;
        RECT 116.310 104.205 117.890 104.535 ;
        RECT 138.505 104.205 140.085 104.535 ;
        RECT 33.510 101.610 34.470 101.760 ;
        RECT 33.510 101.460 47.000 101.610 ;
        RECT 60.825 101.485 62.405 101.815 ;
        RECT 83.020 101.485 84.600 101.815 ;
        RECT 105.215 101.485 106.795 101.815 ;
        RECT 127.410 101.485 128.990 101.815 ;
        RECT 48.745 101.460 49.075 101.475 ;
        RECT 33.510 101.160 49.075 101.460 ;
        RECT 33.510 101.010 47.000 101.160 ;
        RECT 48.745 101.145 49.075 101.160 ;
        RECT 33.510 100.860 34.470 101.010 ;
        RECT 71.920 98.765 73.500 99.095 ;
        RECT 94.115 98.765 95.695 99.095 ;
        RECT 116.310 98.765 117.890 99.095 ;
        RECT 138.505 98.765 140.085 99.095 ;
        RECT 39.530 98.210 40.490 98.360 ;
        RECT 39.530 98.060 47.000 98.210 ;
        RECT 58.865 98.060 59.195 98.075 ;
        RECT 39.530 97.760 59.195 98.060 ;
        RECT 39.530 97.610 47.000 97.760 ;
        RECT 58.865 97.745 59.195 97.760 ;
        RECT 39.530 97.460 40.490 97.610 ;
        RECT 60.825 96.045 62.405 96.375 ;
        RECT 83.020 96.045 84.600 96.375 ;
        RECT 105.215 96.045 106.795 96.375 ;
        RECT 127.410 96.045 128.990 96.375 ;
        RECT 71.920 93.325 73.500 93.655 ;
        RECT 94.115 93.325 95.695 93.655 ;
        RECT 116.310 93.325 117.890 93.655 ;
        RECT 138.505 93.325 140.085 93.655 ;
        RECT 60.825 90.605 62.405 90.935 ;
        RECT 83.020 90.605 84.600 90.935 ;
        RECT 105.215 90.605 106.795 90.935 ;
        RECT 127.410 90.605 128.990 90.935 ;
        RECT 71.920 87.885 73.500 88.215 ;
        RECT 94.115 87.885 95.695 88.215 ;
        RECT 116.310 87.885 117.890 88.215 ;
        RECT 138.505 87.885 140.085 88.215 ;
        RECT 60.825 85.165 62.405 85.495 ;
        RECT 83.020 85.165 84.600 85.495 ;
        RECT 105.215 85.165 106.795 85.495 ;
        RECT 127.410 85.165 128.990 85.495 ;
        RECT 71.920 82.445 73.500 82.775 ;
        RECT 94.115 82.445 95.695 82.775 ;
        RECT 116.310 82.445 117.890 82.775 ;
        RECT 138.505 82.445 140.085 82.775 ;
        RECT 60.825 79.725 62.405 80.055 ;
        RECT 83.020 79.725 84.600 80.055 ;
        RECT 105.215 79.725 106.795 80.055 ;
        RECT 127.410 79.725 128.990 80.055 ;
        RECT 71.920 77.005 73.500 77.335 ;
        RECT 94.115 77.005 95.695 77.335 ;
        RECT 116.310 77.005 117.890 77.335 ;
        RECT 138.505 77.005 140.085 77.335 ;
        RECT 60.825 74.285 62.405 74.615 ;
        RECT 83.020 74.285 84.600 74.615 ;
        RECT 105.215 74.285 106.795 74.615 ;
        RECT 127.410 74.285 128.990 74.615 ;
        RECT 71.920 71.565 73.500 71.895 ;
        RECT 94.115 71.565 95.695 71.895 ;
        RECT 116.310 71.565 117.890 71.895 ;
        RECT 138.505 71.565 140.085 71.895 ;
        RECT 60.825 68.845 62.405 69.175 ;
        RECT 83.020 68.845 84.600 69.175 ;
        RECT 105.215 68.845 106.795 69.175 ;
        RECT 127.410 68.845 128.990 69.175 ;
        RECT 71.920 66.125 73.500 66.455 ;
        RECT 94.115 66.125 95.695 66.455 ;
        RECT 116.310 66.125 117.890 66.455 ;
        RECT 138.505 66.125 140.085 66.455 ;
        RECT 60.825 63.405 62.405 63.735 ;
        RECT 83.020 63.405 84.600 63.735 ;
        RECT 105.215 63.405 106.795 63.735 ;
        RECT 127.410 63.405 128.990 63.735 ;
        RECT 71.920 60.685 73.500 61.015 ;
        RECT 94.115 60.685 95.695 61.015 ;
        RECT 116.310 60.685 117.890 61.015 ;
        RECT 138.505 60.685 140.085 61.015 ;
      LAYER via3 ;
        RECT 71.950 136.850 72.270 137.170 ;
        RECT 72.350 136.850 72.670 137.170 ;
        RECT 72.750 136.850 73.070 137.170 ;
        RECT 73.150 136.850 73.470 137.170 ;
        RECT 94.145 136.850 94.465 137.170 ;
        RECT 94.545 136.850 94.865 137.170 ;
        RECT 94.945 136.850 95.265 137.170 ;
        RECT 95.345 136.850 95.665 137.170 ;
        RECT 116.340 136.850 116.660 137.170 ;
        RECT 116.740 136.850 117.060 137.170 ;
        RECT 117.140 136.850 117.460 137.170 ;
        RECT 117.540 136.850 117.860 137.170 ;
        RECT 138.535 136.850 138.855 137.170 ;
        RECT 138.935 136.850 139.255 137.170 ;
        RECT 139.335 136.850 139.655 137.170 ;
        RECT 139.735 136.850 140.055 137.170 ;
        RECT 60.855 134.130 61.175 134.450 ;
        RECT 61.255 134.130 61.575 134.450 ;
        RECT 61.655 134.130 61.975 134.450 ;
        RECT 62.055 134.130 62.375 134.450 ;
        RECT 83.050 134.130 83.370 134.450 ;
        RECT 83.450 134.130 83.770 134.450 ;
        RECT 83.850 134.130 84.170 134.450 ;
        RECT 84.250 134.130 84.570 134.450 ;
        RECT 105.245 134.130 105.565 134.450 ;
        RECT 105.645 134.130 105.965 134.450 ;
        RECT 106.045 134.130 106.365 134.450 ;
        RECT 106.445 134.130 106.765 134.450 ;
        RECT 127.440 134.130 127.760 134.450 ;
        RECT 127.840 134.130 128.160 134.450 ;
        RECT 128.240 134.130 128.560 134.450 ;
        RECT 128.640 134.130 128.960 134.450 ;
        RECT 71.950 131.410 72.270 131.730 ;
        RECT 72.350 131.410 72.670 131.730 ;
        RECT 72.750 131.410 73.070 131.730 ;
        RECT 73.150 131.410 73.470 131.730 ;
        RECT 94.145 131.410 94.465 131.730 ;
        RECT 94.545 131.410 94.865 131.730 ;
        RECT 94.945 131.410 95.265 131.730 ;
        RECT 95.345 131.410 95.665 131.730 ;
        RECT 116.340 131.410 116.660 131.730 ;
        RECT 116.740 131.410 117.060 131.730 ;
        RECT 117.140 131.410 117.460 131.730 ;
        RECT 117.540 131.410 117.860 131.730 ;
        RECT 138.535 131.410 138.855 131.730 ;
        RECT 138.935 131.410 139.255 131.730 ;
        RECT 139.335 131.410 139.655 131.730 ;
        RECT 139.735 131.410 140.055 131.730 ;
        RECT 60.855 128.690 61.175 129.010 ;
        RECT 61.255 128.690 61.575 129.010 ;
        RECT 61.655 128.690 61.975 129.010 ;
        RECT 62.055 128.690 62.375 129.010 ;
        RECT 83.050 128.690 83.370 129.010 ;
        RECT 83.450 128.690 83.770 129.010 ;
        RECT 83.850 128.690 84.170 129.010 ;
        RECT 84.250 128.690 84.570 129.010 ;
        RECT 105.245 128.690 105.565 129.010 ;
        RECT 105.645 128.690 105.965 129.010 ;
        RECT 106.045 128.690 106.365 129.010 ;
        RECT 106.445 128.690 106.765 129.010 ;
        RECT 127.440 128.690 127.760 129.010 ;
        RECT 127.840 128.690 128.160 129.010 ;
        RECT 128.240 128.690 128.560 129.010 ;
        RECT 128.640 128.690 128.960 129.010 ;
        RECT 71.950 125.970 72.270 126.290 ;
        RECT 72.350 125.970 72.670 126.290 ;
        RECT 72.750 125.970 73.070 126.290 ;
        RECT 73.150 125.970 73.470 126.290 ;
        RECT 94.145 125.970 94.465 126.290 ;
        RECT 94.545 125.970 94.865 126.290 ;
        RECT 94.945 125.970 95.265 126.290 ;
        RECT 95.345 125.970 95.665 126.290 ;
        RECT 116.340 125.970 116.660 126.290 ;
        RECT 116.740 125.970 117.060 126.290 ;
        RECT 117.140 125.970 117.460 126.290 ;
        RECT 117.540 125.970 117.860 126.290 ;
        RECT 138.535 125.970 138.855 126.290 ;
        RECT 138.935 125.970 139.255 126.290 ;
        RECT 139.335 125.970 139.655 126.290 ;
        RECT 139.735 125.970 140.055 126.290 ;
        RECT 60.855 123.250 61.175 123.570 ;
        RECT 61.255 123.250 61.575 123.570 ;
        RECT 61.655 123.250 61.975 123.570 ;
        RECT 62.055 123.250 62.375 123.570 ;
        RECT 83.050 123.250 83.370 123.570 ;
        RECT 83.450 123.250 83.770 123.570 ;
        RECT 83.850 123.250 84.170 123.570 ;
        RECT 84.250 123.250 84.570 123.570 ;
        RECT 105.245 123.250 105.565 123.570 ;
        RECT 105.645 123.250 105.965 123.570 ;
        RECT 106.045 123.250 106.365 123.570 ;
        RECT 106.445 123.250 106.765 123.570 ;
        RECT 127.440 123.250 127.760 123.570 ;
        RECT 127.840 123.250 128.160 123.570 ;
        RECT 128.240 123.250 128.560 123.570 ;
        RECT 128.640 123.250 128.960 123.570 ;
        RECT 71.950 120.530 72.270 120.850 ;
        RECT 72.350 120.530 72.670 120.850 ;
        RECT 72.750 120.530 73.070 120.850 ;
        RECT 73.150 120.530 73.470 120.850 ;
        RECT 94.145 120.530 94.465 120.850 ;
        RECT 94.545 120.530 94.865 120.850 ;
        RECT 94.945 120.530 95.265 120.850 ;
        RECT 95.345 120.530 95.665 120.850 ;
        RECT 116.340 120.530 116.660 120.850 ;
        RECT 116.740 120.530 117.060 120.850 ;
        RECT 117.140 120.530 117.460 120.850 ;
        RECT 117.540 120.530 117.860 120.850 ;
        RECT 138.535 120.530 138.855 120.850 ;
        RECT 138.935 120.530 139.255 120.850 ;
        RECT 139.335 120.530 139.655 120.850 ;
        RECT 139.735 120.530 140.055 120.850 ;
        RECT 60.855 117.810 61.175 118.130 ;
        RECT 61.255 117.810 61.575 118.130 ;
        RECT 61.655 117.810 61.975 118.130 ;
        RECT 62.055 117.810 62.375 118.130 ;
        RECT 83.050 117.810 83.370 118.130 ;
        RECT 83.450 117.810 83.770 118.130 ;
        RECT 83.850 117.810 84.170 118.130 ;
        RECT 84.250 117.810 84.570 118.130 ;
        RECT 105.245 117.810 105.565 118.130 ;
        RECT 105.645 117.810 105.965 118.130 ;
        RECT 106.045 117.810 106.365 118.130 ;
        RECT 106.445 117.810 106.765 118.130 ;
        RECT 127.440 117.810 127.760 118.130 ;
        RECT 127.840 117.810 128.160 118.130 ;
        RECT 128.240 117.810 128.560 118.130 ;
        RECT 128.640 117.810 128.960 118.130 ;
        RECT 71.950 115.090 72.270 115.410 ;
        RECT 72.350 115.090 72.670 115.410 ;
        RECT 72.750 115.090 73.070 115.410 ;
        RECT 73.150 115.090 73.470 115.410 ;
        RECT 94.145 115.090 94.465 115.410 ;
        RECT 94.545 115.090 94.865 115.410 ;
        RECT 94.945 115.090 95.265 115.410 ;
        RECT 95.345 115.090 95.665 115.410 ;
        RECT 116.340 115.090 116.660 115.410 ;
        RECT 116.740 115.090 117.060 115.410 ;
        RECT 117.140 115.090 117.460 115.410 ;
        RECT 117.540 115.090 117.860 115.410 ;
        RECT 138.535 115.090 138.855 115.410 ;
        RECT 138.935 115.090 139.255 115.410 ;
        RECT 139.335 115.090 139.655 115.410 ;
        RECT 139.735 115.090 140.055 115.410 ;
        RECT 60.855 112.370 61.175 112.690 ;
        RECT 61.255 112.370 61.575 112.690 ;
        RECT 61.655 112.370 61.975 112.690 ;
        RECT 62.055 112.370 62.375 112.690 ;
        RECT 83.050 112.370 83.370 112.690 ;
        RECT 83.450 112.370 83.770 112.690 ;
        RECT 83.850 112.370 84.170 112.690 ;
        RECT 84.250 112.370 84.570 112.690 ;
        RECT 105.245 112.370 105.565 112.690 ;
        RECT 105.645 112.370 105.965 112.690 ;
        RECT 106.045 112.370 106.365 112.690 ;
        RECT 106.445 112.370 106.765 112.690 ;
        RECT 127.440 112.370 127.760 112.690 ;
        RECT 127.840 112.370 128.160 112.690 ;
        RECT 128.240 112.370 128.560 112.690 ;
        RECT 128.640 112.370 128.960 112.690 ;
        RECT 71.950 109.650 72.270 109.970 ;
        RECT 72.350 109.650 72.670 109.970 ;
        RECT 72.750 109.650 73.070 109.970 ;
        RECT 73.150 109.650 73.470 109.970 ;
        RECT 94.145 109.650 94.465 109.970 ;
        RECT 94.545 109.650 94.865 109.970 ;
        RECT 94.945 109.650 95.265 109.970 ;
        RECT 95.345 109.650 95.665 109.970 ;
        RECT 116.340 109.650 116.660 109.970 ;
        RECT 116.740 109.650 117.060 109.970 ;
        RECT 117.140 109.650 117.460 109.970 ;
        RECT 117.540 109.650 117.860 109.970 ;
        RECT 138.535 109.650 138.855 109.970 ;
        RECT 138.935 109.650 139.255 109.970 ;
        RECT 139.335 109.650 139.655 109.970 ;
        RECT 139.735 109.650 140.055 109.970 ;
        RECT 60.855 106.930 61.175 107.250 ;
        RECT 61.255 106.930 61.575 107.250 ;
        RECT 61.655 106.930 61.975 107.250 ;
        RECT 62.055 106.930 62.375 107.250 ;
        RECT 83.050 106.930 83.370 107.250 ;
        RECT 83.450 106.930 83.770 107.250 ;
        RECT 83.850 106.930 84.170 107.250 ;
        RECT 84.250 106.930 84.570 107.250 ;
        RECT 105.245 106.930 105.565 107.250 ;
        RECT 105.645 106.930 105.965 107.250 ;
        RECT 106.045 106.930 106.365 107.250 ;
        RECT 106.445 106.930 106.765 107.250 ;
        RECT 127.440 106.930 127.760 107.250 ;
        RECT 127.840 106.930 128.160 107.250 ;
        RECT 128.240 106.930 128.560 107.250 ;
        RECT 128.640 106.930 128.960 107.250 ;
        RECT 37.250 104.350 37.970 105.070 ;
        RECT 71.950 104.210 72.270 104.530 ;
        RECT 72.350 104.210 72.670 104.530 ;
        RECT 72.750 104.210 73.070 104.530 ;
        RECT 73.150 104.210 73.470 104.530 ;
        RECT 94.145 104.210 94.465 104.530 ;
        RECT 94.545 104.210 94.865 104.530 ;
        RECT 94.945 104.210 95.265 104.530 ;
        RECT 95.345 104.210 95.665 104.530 ;
        RECT 116.340 104.210 116.660 104.530 ;
        RECT 116.740 104.210 117.060 104.530 ;
        RECT 117.140 104.210 117.460 104.530 ;
        RECT 117.540 104.210 117.860 104.530 ;
        RECT 138.535 104.210 138.855 104.530 ;
        RECT 138.935 104.210 139.255 104.530 ;
        RECT 139.335 104.210 139.655 104.530 ;
        RECT 139.735 104.210 140.055 104.530 ;
        RECT 33.630 100.950 34.350 101.670 ;
        RECT 60.855 101.490 61.175 101.810 ;
        RECT 61.255 101.490 61.575 101.810 ;
        RECT 61.655 101.490 61.975 101.810 ;
        RECT 62.055 101.490 62.375 101.810 ;
        RECT 83.050 101.490 83.370 101.810 ;
        RECT 83.450 101.490 83.770 101.810 ;
        RECT 83.850 101.490 84.170 101.810 ;
        RECT 84.250 101.490 84.570 101.810 ;
        RECT 105.245 101.490 105.565 101.810 ;
        RECT 105.645 101.490 105.965 101.810 ;
        RECT 106.045 101.490 106.365 101.810 ;
        RECT 106.445 101.490 106.765 101.810 ;
        RECT 127.440 101.490 127.760 101.810 ;
        RECT 127.840 101.490 128.160 101.810 ;
        RECT 128.240 101.490 128.560 101.810 ;
        RECT 128.640 101.490 128.960 101.810 ;
        RECT 71.950 98.770 72.270 99.090 ;
        RECT 72.350 98.770 72.670 99.090 ;
        RECT 72.750 98.770 73.070 99.090 ;
        RECT 73.150 98.770 73.470 99.090 ;
        RECT 94.145 98.770 94.465 99.090 ;
        RECT 94.545 98.770 94.865 99.090 ;
        RECT 94.945 98.770 95.265 99.090 ;
        RECT 95.345 98.770 95.665 99.090 ;
        RECT 116.340 98.770 116.660 99.090 ;
        RECT 116.740 98.770 117.060 99.090 ;
        RECT 117.140 98.770 117.460 99.090 ;
        RECT 117.540 98.770 117.860 99.090 ;
        RECT 138.535 98.770 138.855 99.090 ;
        RECT 138.935 98.770 139.255 99.090 ;
        RECT 139.335 98.770 139.655 99.090 ;
        RECT 139.735 98.770 140.055 99.090 ;
        RECT 39.650 97.550 40.370 98.270 ;
        RECT 60.855 96.050 61.175 96.370 ;
        RECT 61.255 96.050 61.575 96.370 ;
        RECT 61.655 96.050 61.975 96.370 ;
        RECT 62.055 96.050 62.375 96.370 ;
        RECT 83.050 96.050 83.370 96.370 ;
        RECT 83.450 96.050 83.770 96.370 ;
        RECT 83.850 96.050 84.170 96.370 ;
        RECT 84.250 96.050 84.570 96.370 ;
        RECT 105.245 96.050 105.565 96.370 ;
        RECT 105.645 96.050 105.965 96.370 ;
        RECT 106.045 96.050 106.365 96.370 ;
        RECT 106.445 96.050 106.765 96.370 ;
        RECT 127.440 96.050 127.760 96.370 ;
        RECT 127.840 96.050 128.160 96.370 ;
        RECT 128.240 96.050 128.560 96.370 ;
        RECT 128.640 96.050 128.960 96.370 ;
        RECT 71.950 93.330 72.270 93.650 ;
        RECT 72.350 93.330 72.670 93.650 ;
        RECT 72.750 93.330 73.070 93.650 ;
        RECT 73.150 93.330 73.470 93.650 ;
        RECT 94.145 93.330 94.465 93.650 ;
        RECT 94.545 93.330 94.865 93.650 ;
        RECT 94.945 93.330 95.265 93.650 ;
        RECT 95.345 93.330 95.665 93.650 ;
        RECT 116.340 93.330 116.660 93.650 ;
        RECT 116.740 93.330 117.060 93.650 ;
        RECT 117.140 93.330 117.460 93.650 ;
        RECT 117.540 93.330 117.860 93.650 ;
        RECT 138.535 93.330 138.855 93.650 ;
        RECT 138.935 93.330 139.255 93.650 ;
        RECT 139.335 93.330 139.655 93.650 ;
        RECT 139.735 93.330 140.055 93.650 ;
        RECT 60.855 90.610 61.175 90.930 ;
        RECT 61.255 90.610 61.575 90.930 ;
        RECT 61.655 90.610 61.975 90.930 ;
        RECT 62.055 90.610 62.375 90.930 ;
        RECT 83.050 90.610 83.370 90.930 ;
        RECT 83.450 90.610 83.770 90.930 ;
        RECT 83.850 90.610 84.170 90.930 ;
        RECT 84.250 90.610 84.570 90.930 ;
        RECT 105.245 90.610 105.565 90.930 ;
        RECT 105.645 90.610 105.965 90.930 ;
        RECT 106.045 90.610 106.365 90.930 ;
        RECT 106.445 90.610 106.765 90.930 ;
        RECT 127.440 90.610 127.760 90.930 ;
        RECT 127.840 90.610 128.160 90.930 ;
        RECT 128.240 90.610 128.560 90.930 ;
        RECT 128.640 90.610 128.960 90.930 ;
        RECT 71.950 87.890 72.270 88.210 ;
        RECT 72.350 87.890 72.670 88.210 ;
        RECT 72.750 87.890 73.070 88.210 ;
        RECT 73.150 87.890 73.470 88.210 ;
        RECT 94.145 87.890 94.465 88.210 ;
        RECT 94.545 87.890 94.865 88.210 ;
        RECT 94.945 87.890 95.265 88.210 ;
        RECT 95.345 87.890 95.665 88.210 ;
        RECT 116.340 87.890 116.660 88.210 ;
        RECT 116.740 87.890 117.060 88.210 ;
        RECT 117.140 87.890 117.460 88.210 ;
        RECT 117.540 87.890 117.860 88.210 ;
        RECT 138.535 87.890 138.855 88.210 ;
        RECT 138.935 87.890 139.255 88.210 ;
        RECT 139.335 87.890 139.655 88.210 ;
        RECT 139.735 87.890 140.055 88.210 ;
        RECT 60.855 85.170 61.175 85.490 ;
        RECT 61.255 85.170 61.575 85.490 ;
        RECT 61.655 85.170 61.975 85.490 ;
        RECT 62.055 85.170 62.375 85.490 ;
        RECT 83.050 85.170 83.370 85.490 ;
        RECT 83.450 85.170 83.770 85.490 ;
        RECT 83.850 85.170 84.170 85.490 ;
        RECT 84.250 85.170 84.570 85.490 ;
        RECT 105.245 85.170 105.565 85.490 ;
        RECT 105.645 85.170 105.965 85.490 ;
        RECT 106.045 85.170 106.365 85.490 ;
        RECT 106.445 85.170 106.765 85.490 ;
        RECT 127.440 85.170 127.760 85.490 ;
        RECT 127.840 85.170 128.160 85.490 ;
        RECT 128.240 85.170 128.560 85.490 ;
        RECT 128.640 85.170 128.960 85.490 ;
        RECT 71.950 82.450 72.270 82.770 ;
        RECT 72.350 82.450 72.670 82.770 ;
        RECT 72.750 82.450 73.070 82.770 ;
        RECT 73.150 82.450 73.470 82.770 ;
        RECT 94.145 82.450 94.465 82.770 ;
        RECT 94.545 82.450 94.865 82.770 ;
        RECT 94.945 82.450 95.265 82.770 ;
        RECT 95.345 82.450 95.665 82.770 ;
        RECT 116.340 82.450 116.660 82.770 ;
        RECT 116.740 82.450 117.060 82.770 ;
        RECT 117.140 82.450 117.460 82.770 ;
        RECT 117.540 82.450 117.860 82.770 ;
        RECT 138.535 82.450 138.855 82.770 ;
        RECT 138.935 82.450 139.255 82.770 ;
        RECT 139.335 82.450 139.655 82.770 ;
        RECT 139.735 82.450 140.055 82.770 ;
        RECT 60.855 79.730 61.175 80.050 ;
        RECT 61.255 79.730 61.575 80.050 ;
        RECT 61.655 79.730 61.975 80.050 ;
        RECT 62.055 79.730 62.375 80.050 ;
        RECT 83.050 79.730 83.370 80.050 ;
        RECT 83.450 79.730 83.770 80.050 ;
        RECT 83.850 79.730 84.170 80.050 ;
        RECT 84.250 79.730 84.570 80.050 ;
        RECT 105.245 79.730 105.565 80.050 ;
        RECT 105.645 79.730 105.965 80.050 ;
        RECT 106.045 79.730 106.365 80.050 ;
        RECT 106.445 79.730 106.765 80.050 ;
        RECT 127.440 79.730 127.760 80.050 ;
        RECT 127.840 79.730 128.160 80.050 ;
        RECT 128.240 79.730 128.560 80.050 ;
        RECT 128.640 79.730 128.960 80.050 ;
        RECT 71.950 77.010 72.270 77.330 ;
        RECT 72.350 77.010 72.670 77.330 ;
        RECT 72.750 77.010 73.070 77.330 ;
        RECT 73.150 77.010 73.470 77.330 ;
        RECT 94.145 77.010 94.465 77.330 ;
        RECT 94.545 77.010 94.865 77.330 ;
        RECT 94.945 77.010 95.265 77.330 ;
        RECT 95.345 77.010 95.665 77.330 ;
        RECT 116.340 77.010 116.660 77.330 ;
        RECT 116.740 77.010 117.060 77.330 ;
        RECT 117.140 77.010 117.460 77.330 ;
        RECT 117.540 77.010 117.860 77.330 ;
        RECT 138.535 77.010 138.855 77.330 ;
        RECT 138.935 77.010 139.255 77.330 ;
        RECT 139.335 77.010 139.655 77.330 ;
        RECT 139.735 77.010 140.055 77.330 ;
        RECT 60.855 74.290 61.175 74.610 ;
        RECT 61.255 74.290 61.575 74.610 ;
        RECT 61.655 74.290 61.975 74.610 ;
        RECT 62.055 74.290 62.375 74.610 ;
        RECT 83.050 74.290 83.370 74.610 ;
        RECT 83.450 74.290 83.770 74.610 ;
        RECT 83.850 74.290 84.170 74.610 ;
        RECT 84.250 74.290 84.570 74.610 ;
        RECT 105.245 74.290 105.565 74.610 ;
        RECT 105.645 74.290 105.965 74.610 ;
        RECT 106.045 74.290 106.365 74.610 ;
        RECT 106.445 74.290 106.765 74.610 ;
        RECT 127.440 74.290 127.760 74.610 ;
        RECT 127.840 74.290 128.160 74.610 ;
        RECT 128.240 74.290 128.560 74.610 ;
        RECT 128.640 74.290 128.960 74.610 ;
        RECT 71.950 71.570 72.270 71.890 ;
        RECT 72.350 71.570 72.670 71.890 ;
        RECT 72.750 71.570 73.070 71.890 ;
        RECT 73.150 71.570 73.470 71.890 ;
        RECT 94.145 71.570 94.465 71.890 ;
        RECT 94.545 71.570 94.865 71.890 ;
        RECT 94.945 71.570 95.265 71.890 ;
        RECT 95.345 71.570 95.665 71.890 ;
        RECT 116.340 71.570 116.660 71.890 ;
        RECT 116.740 71.570 117.060 71.890 ;
        RECT 117.140 71.570 117.460 71.890 ;
        RECT 117.540 71.570 117.860 71.890 ;
        RECT 138.535 71.570 138.855 71.890 ;
        RECT 138.935 71.570 139.255 71.890 ;
        RECT 139.335 71.570 139.655 71.890 ;
        RECT 139.735 71.570 140.055 71.890 ;
        RECT 60.855 68.850 61.175 69.170 ;
        RECT 61.255 68.850 61.575 69.170 ;
        RECT 61.655 68.850 61.975 69.170 ;
        RECT 62.055 68.850 62.375 69.170 ;
        RECT 83.050 68.850 83.370 69.170 ;
        RECT 83.450 68.850 83.770 69.170 ;
        RECT 83.850 68.850 84.170 69.170 ;
        RECT 84.250 68.850 84.570 69.170 ;
        RECT 105.245 68.850 105.565 69.170 ;
        RECT 105.645 68.850 105.965 69.170 ;
        RECT 106.045 68.850 106.365 69.170 ;
        RECT 106.445 68.850 106.765 69.170 ;
        RECT 127.440 68.850 127.760 69.170 ;
        RECT 127.840 68.850 128.160 69.170 ;
        RECT 128.240 68.850 128.560 69.170 ;
        RECT 128.640 68.850 128.960 69.170 ;
        RECT 71.950 66.130 72.270 66.450 ;
        RECT 72.350 66.130 72.670 66.450 ;
        RECT 72.750 66.130 73.070 66.450 ;
        RECT 73.150 66.130 73.470 66.450 ;
        RECT 94.145 66.130 94.465 66.450 ;
        RECT 94.545 66.130 94.865 66.450 ;
        RECT 94.945 66.130 95.265 66.450 ;
        RECT 95.345 66.130 95.665 66.450 ;
        RECT 116.340 66.130 116.660 66.450 ;
        RECT 116.740 66.130 117.060 66.450 ;
        RECT 117.140 66.130 117.460 66.450 ;
        RECT 117.540 66.130 117.860 66.450 ;
        RECT 138.535 66.130 138.855 66.450 ;
        RECT 138.935 66.130 139.255 66.450 ;
        RECT 139.335 66.130 139.655 66.450 ;
        RECT 139.735 66.130 140.055 66.450 ;
        RECT 60.855 63.410 61.175 63.730 ;
        RECT 61.255 63.410 61.575 63.730 ;
        RECT 61.655 63.410 61.975 63.730 ;
        RECT 62.055 63.410 62.375 63.730 ;
        RECT 83.050 63.410 83.370 63.730 ;
        RECT 83.450 63.410 83.770 63.730 ;
        RECT 83.850 63.410 84.170 63.730 ;
        RECT 84.250 63.410 84.570 63.730 ;
        RECT 105.245 63.410 105.565 63.730 ;
        RECT 105.645 63.410 105.965 63.730 ;
        RECT 106.045 63.410 106.365 63.730 ;
        RECT 106.445 63.410 106.765 63.730 ;
        RECT 127.440 63.410 127.760 63.730 ;
        RECT 127.840 63.410 128.160 63.730 ;
        RECT 128.240 63.410 128.560 63.730 ;
        RECT 128.640 63.410 128.960 63.730 ;
        RECT 71.950 60.690 72.270 61.010 ;
        RECT 72.350 60.690 72.670 61.010 ;
        RECT 72.750 60.690 73.070 61.010 ;
        RECT 73.150 60.690 73.470 61.010 ;
        RECT 94.145 60.690 94.465 61.010 ;
        RECT 94.545 60.690 94.865 61.010 ;
        RECT 94.945 60.690 95.265 61.010 ;
        RECT 95.345 60.690 95.665 61.010 ;
        RECT 116.340 60.690 116.660 61.010 ;
        RECT 116.740 60.690 117.060 61.010 ;
        RECT 117.140 60.690 117.460 61.010 ;
        RECT 117.540 60.690 117.860 61.010 ;
        RECT 138.535 60.690 138.855 61.010 ;
        RECT 138.935 60.690 139.255 61.010 ;
        RECT 139.335 60.690 139.655 61.010 ;
        RECT 139.735 60.690 140.055 61.010 ;
      LAYER met4 ;
        RECT 6.000 4.970 8.000 220.730 ;
        RECT 9.000 220.440 11.000 220.730 ;
        RECT 35.670 220.440 35.970 225.730 ;
        RECT 38.430 220.440 38.730 225.730 ;
        RECT 41.190 220.440 41.490 225.730 ;
        RECT 43.950 220.440 44.250 225.730 ;
        RECT 46.710 220.440 47.010 225.730 ;
        RECT 49.470 220.440 49.770 225.730 ;
        RECT 52.230 220.440 52.530 225.730 ;
        RECT 54.990 220.440 55.290 225.730 ;
        RECT 57.750 220.440 58.050 225.730 ;
        RECT 60.510 220.440 60.810 225.730 ;
        RECT 63.270 220.440 63.570 225.730 ;
        RECT 66.030 220.440 66.330 225.730 ;
        RECT 68.790 220.440 69.090 225.730 ;
        RECT 71.550 220.440 71.850 225.730 ;
        RECT 74.310 220.440 74.610 225.730 ;
        RECT 77.070 220.440 77.370 225.730 ;
        RECT 79.830 224.730 80.130 225.730 ;
        RECT 82.590 224.730 82.890 225.730 ;
        RECT 85.350 224.730 85.650 225.730 ;
        RECT 88.110 224.730 88.410 225.730 ;
        RECT 90.870 224.730 91.170 225.730 ;
        RECT 93.630 224.730 93.930 225.730 ;
        RECT 96.390 224.730 96.690 225.730 ;
        RECT 99.150 224.730 99.450 225.730 ;
        RECT 101.910 224.730 102.210 225.730 ;
        RECT 104.670 224.730 104.970 225.730 ;
        RECT 107.430 224.730 107.730 225.730 ;
        RECT 110.190 224.730 110.490 225.730 ;
        RECT 112.950 224.730 113.250 225.730 ;
        RECT 115.710 224.730 116.010 225.730 ;
        RECT 118.470 224.730 118.770 225.730 ;
        RECT 121.230 224.730 121.530 225.730 ;
        RECT 123.990 224.730 124.290 225.730 ;
        RECT 126.750 224.730 127.050 225.730 ;
        RECT 129.510 224.730 129.810 225.730 ;
        RECT 132.270 224.730 132.570 225.730 ;
        RECT 135.030 224.730 135.330 225.730 ;
        RECT 137.790 224.730 138.090 225.730 ;
        RECT 140.550 224.730 140.850 225.730 ;
        RECT 143.310 224.730 143.610 225.730 ;
        RECT 146.070 224.730 146.370 225.730 ;
        RECT 148.830 224.730 149.130 225.730 ;
        RECT 151.590 224.730 151.890 225.730 ;
        RECT 9.000 218.440 86.820 220.440 ;
        RECT 9.000 4.970 11.000 218.440 ;
        RECT 32.800 161.440 157.710 162.340 ;
        RECT 32.800 105.110 33.700 161.440 ;
        RECT 37.155 105.110 38.065 105.165 ;
        RECT 32.800 104.210 38.720 105.110 ;
        RECT 33.535 101.760 34.445 101.765 ;
        RECT 28.700 100.860 38.660 101.760 ;
        RECT 28.700 42.850 29.600 100.860 ;
        RECT 33.535 100.855 34.445 100.860 ;
        RECT 39.555 98.340 40.465 98.365 ;
        RECT 37.690 97.440 42.110 98.340 ;
        RECT 37.690 51.230 38.590 97.440 ;
        RECT 60.815 60.610 62.415 137.250 ;
        RECT 71.910 60.610 73.510 137.250 ;
        RECT 83.010 60.610 84.610 137.250 ;
        RECT 94.105 60.610 95.705 137.250 ;
        RECT 105.205 60.610 106.805 137.250 ;
        RECT 116.300 60.610 117.900 137.250 ;
        RECT 127.400 60.610 129.000 137.250 ;
        RECT 138.495 60.610 140.095 137.250 ;
        RECT 37.690 50.330 138.390 51.230 ;
        RECT 28.700 41.950 119.070 42.850 ;
        RECT 21.570 -0.030 22.470 0.970 ;
        RECT 40.890 -0.030 41.790 0.970 ;
        RECT 60.210 -0.030 61.110 0.970 ;
        RECT 79.530 -0.030 80.430 0.970 ;
        RECT 98.850 -0.030 99.750 0.970 ;
        RECT 118.170 -0.030 119.070 41.950 ;
        RECT 137.490 -0.030 138.390 50.330 ;
        RECT 156.810 -0.030 157.710 161.440 ;
  END
END tt_um_brandonramos_opamp_ladder
END LIBRARY

